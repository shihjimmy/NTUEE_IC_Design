`timescale 1ns/1ps
`define SIZE 10000
module tb_kendall();

	wire [3:0] i0_x, i1_x, i2_x, i3_x;
	wire [3:0] i0_y, i1_y, i2_y, i3_y;
	wire [3:0] kendall;

	reg  [3:0] i0mem[0:2*`SIZE-1];
	reg  [3:0] i1mem[0:2*`SIZE-1];
	reg  [3:0] i2mem[0:2*`SIZE-1];
	reg  [3:0] i3mem[0:2*`SIZE-1];

	reg  [3:0] kendallmem[0:`SIZE-1];
	wire  [3:0] ans;


	integer i,j,error,error_total,error_part,hide;
	integer err3,err4,err5,err6, err7,err10,err20;
	real time_avg,time_step_sum,time_step,acc,total;




	kendall_rank top(					.kendall(kendall),
										.i0_x(i0_x),
										.i0_y(i0_y),
										.i1_x(i1_x),
										.i1_y(i1_y),
										.i2_x(i2_x),
										.i2_y(i2_y),
										.i3_x(i3_x),
										.i3_y(i3_y)
										);


	initial	begin
		$readmemh("i0.dat", i0mem);
		$readmemh("i1.dat", i1mem);
		$readmemh("i2.dat", i2mem);
		$readmemh("i3.dat", i3mem);
		$readmemb("golden.dat",kendallmem);


	end
	initial begin
		$fsdbDumpfile("kendall.fsdb");
		$fsdbDumpvars;
		$fsdbDumpMDA;
	end

	initial
	begin
		i = 0;
		err3 = 0;
		err4 = 0;
		err5 = 0;
		err6 = 0;
		err7 = 0;
		err10 = 0;
		err20 = 0;
	end

	assign i0_x  = i0mem[i];
	assign i0_y  = i0mem[i+1];
	assign i1_x  = i1mem[i];
	assign i1_y  = i1mem[i+1];
	assign i2_x  = i2mem[i];
	assign i2_y  = i2mem[i+1];
	assign i3_x  = i3mem[i];
	assign i3_y  = i3mem[i+1];

	assign ans = kendallmem[i/2];

	always begin
		#3.5
		if(ans!==kendall)
			err3 = err3 + 1;
	    #0.5
		if(ans!==kendall)
			err4 = err4 + 1;
		#0.5
		if(ans!==kendall)
			err5 = err5 + 1;
		#0.5
		if(ans!==kendall)
			err6 = err6 + 1;
		#0.5
		if(ans!==kendall)
			err7 = err7 + 1;
		#0.5
		if(ans!==kendall)
			err10 = err10 + 1;
		#14
		if(ans!==kendall)
			err20 = err20 + 1;
		#1
		i = i + 2;
	end

	always @(i) begin
		if(i == 10000) begin
		    if(err3 == 0) begin
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;130m▒\033[38;5;214;48;5;137m▒\033[38;5;178;48;5;188m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;130;48;5;187m▒\033[38;5;130;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;180;48;5;224m░\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;179m▒\033[38;5;178;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;230m░\033[38;5;214;48;5;143m▒\033[38;5;172;48;5;136m▒\033[38;5;130;48;5;216m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;137;48;5;187m▒\033[38;5;221;48;5;101m▒\033[38;5;172;48;5;58m░\033[38;5;208;48;5;52m░\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;130m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;180m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;187m▒\033[38;5;221;48;5;101m▒\033[38;5;172;48;5;95m▒\033[38;5;215;48;5;52m \033[38;5;172;48;5;58m░\033[38;5;172;48;5;136m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;180m▒\033[38;5;214;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;179;48;5;223m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;94m░\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;172;48;5;216m░\033[38;5;179;48;5;222m░\033[38;5;221;48;5;185m░\033[38;5;136;48;5;185m░\033[38;5;214;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;223;48;5;224m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;172;48;5;137m▒\033[38;5;208;48;5;58m▒\033[38;5;202;48;5;239m▒\033[38;5;166;48;5;137m▓\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;130;48;5;58m▒\033[38;5;173;48;5;238m▓\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;229m \033[38;5;221;48;5;187m▒\033[38;5;94;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m░\033[38;5;214;48;5;186m░\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;58m▒\033[38;5;221;48;5;58m▒\033[38;5;179;48;5;58m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;221m░\033[38;5;214;48;5;221m░\033[38;5;94;48;5;185m░\033[38;5;136;48;5;186m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;185m▒\033[38;5;220;48;5;222m░\033[38;5;229;48;5;229m \033[38;5;221;48;5;224m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;130;48;5;230m \033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;222m░\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;230m \033[38;5;221;48;5;230m░\033[38;5;221;48;5;230m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;221;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;180m▓\033[38;5;166;48;5;235m▒\033[38;5;16;48;5;16m▓\033[38;5;216;48;5;232m░\033[38;5;173;48;5;233m▒\033[38;5;94;48;5;144m▓\033[38;5;220;48;5;223m▒\033[38;5;185;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;220;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;144m▓\033[38;5;179;48;5;138m▓\033[38;5;172;48;5;95m▓\033[38;5;130;48;5;236m▓\033[38;5;173;48;5;235m▓\033[38;5;166;48;5;236m▓\033[38;5;94;48;5;101m▓\033[38;5;220;48;5;187m▒\033[38;5;185;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;136;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;143m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;58m▒\033[38;5;214;48;5;58m▒\033[38;5;221;48;5;234m░\033[38;5;178;48;5;234m░\033[38;5;220;48;5;233m \033[38;5;185;48;5;235m▒\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;223m▒\033[38;5;136;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;187m▒\033[38;5;136;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;136;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;136;48;5;223m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;179;48;5;186m░\033[38;5;172;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;214;48;5;223m░\033[38;5;94;48;5;223m░\033[38;5;221;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;202;48;5;224m░\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;178;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;136;48;5;180m▒\033[38;5;172;48;5;187m▒\033[38;5;209;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;220;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;130;48;5;224m░\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;173m▒\033[38;5;214;48;5;173m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;221;48;5;223m░\033[38;5;221;48;5;223m░\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;180m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;187m▒\033[38;5;136;48;5;230m░\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;172;48;5;224m░\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;187m▒\033[38;5;214;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;231m \033[38;5;172;48;5;224m \033[38;5;179;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;214;48;5;223m░\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;186m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;130;48;5;255m░\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;186m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;172;48;5;187m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;214;48;5;187m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;172;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;178;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;230m \033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;186m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;231m \033[38;5;172;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;178;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;223m░\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;136;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;214;48;5;187m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;178;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;230m \033[38;5;179;48;5;186m░\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;230m \033[38;5;136;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;223m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;101m▓\033[38;5;214;48;5;235m▒\033[38;5;94;48;5;234m▒\033[38;5;94;48;5;234m▒\033[38;5;94;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;94;48;5;234m▒\033[38;5;94;48;5;234m▒\033[38;5;94;48;5;234m▒\033[38;5;94;48;5;237m▒\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;95m▓\033[38;5;94;48;5;235m▒\033[38;5;221;48;5;234m▒\033[38;5;221;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;94;48;5;236m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;59m▓\033[38;5;94;48;5;236m▒\033[38;5;179;48;5;234m▒\033[38;5;172;48;5;234m░\033[38;5;172;48;5;235m░\033[38;5;172;48;5;58m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;95m▓\033[38;5;94;48;5;237m▓\033[38;5;179;48;5;234m▒\033[38;5;94;48;5;234m▒\033[38;5;214;48;5;236m▒\033[38;5;214;48;5;240m▓\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;223m░\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;178;48;5;187m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;222;48;5;232m \033[38;5;94;48;5;137m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;233m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;236m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;238m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;186m░\033[38;5;214;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;187m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;250;48;5;249m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;221;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;240;48;5;240m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;237;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;232m \033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;180m▒\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;187m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;137m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;232m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;246;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;239;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;242m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;232;48;5;232m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;243;48;5;242m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;246;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;239;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;179;48;5;94m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;186m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;187m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;235;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;253m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;236;48;5;235m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;232;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;232m \033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;222;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;230m░\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;223m░\033[38;5;178;48;5;230m \033[38;5;179;48;5;186m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;232m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;245;48;5;245m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;248m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;246;48;5;246m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;246;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;178;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;186m░\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;136;48;5;223m░\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;137m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;234;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;237m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;232;48;5;232m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;252m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;179;48;5;234m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;186m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;223m░\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;222;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;137m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;240;48;5;240m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;7;48;5;7m▓\033[38;5;235;48;5;235m▓\033[38;5;232;48;5;232m▓\033[38;5;232;48;5;232m▓\033[38;5;236;48;5;235m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;236;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;145;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;236;48;5;235m▓\033[38;5;232;48;5;232m▓\033[38;5;232;48;5;232m▓\033[38;5;235;48;5;235m▓\033[38;5;7;48;5;7m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;245;48;5;245m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;130;48;5;237m▓\033[38;5;166;48;5;223m░\033[38;5;208;48;5;224m \033[38;5;130;48;5;223m░\033[38;5;208;48;5;180m▒\033[38;5;208;48;5;173m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;136;48;5;144m▓\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;220;48;5;179m▒\033[38;5;178;48;5;229m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;230m \033[38;5;214;48;5;180m▒\033[38;5;94;48;5;137m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;234;48;5;234m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;236m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;233;48;5;233m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;249;48;5;249m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;102;48;5;102m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;252;48;5;252m▓\033[38;5;241;48;5;59m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;243;48;5;243m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;188m▓\033[38;5;243;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;232m░\033[38;5;172;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;130;48;5;230m \033[38;5;130;48;5;223m░\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;187m▒\033[38;5;178;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;214;48;5;186m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;214;48;5;230m░\033[38;5;94;48;5;180m▓\033[38;5;214;48;5;233m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;58m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;235m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;233m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;136;48;5;234m▒\033[38;5;94;48;5;143m▓\033[38;5;179;48;5;187m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;223m░\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;178;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;230m░\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m░\033[38;5;214;48;5;180m░\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;222;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;172;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;130;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;179;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;230m \033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;223m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;229m \033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;216;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;172;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;172;48;5;187m▒\033[38;5;221;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;223m░\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m░\033[38;5;178;48;5;186m░\033[38;5;136;48;5;185m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;178;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;216;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;172;48;5;180m▒\033[38;5;172;48;5;173m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;172;48;5;223m░\033[38;5;209;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;222m░\033[38;5;136;48;5;186m░\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;223m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;202;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;223m░\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;186m░\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;216;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;186m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;172;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;223m░\033[38;5;220;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;187m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;220;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;172;48;5;223m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;179;48;5;223m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;178;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;230m \033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;179;48;5;143m▓\033[38;5;172;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;136;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;221;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;179;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;144m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;137m▓\033[38;5;220;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;136;48;5;186m▒\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;222;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;144m▓\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;178;48;5;179m▒\033[38;5;220;48;5;179m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;178;48;5;186m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;178;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;101m▒\033[38;5;220;48;5;137m▓\033[38;5;230;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;130;48;5;230m \033[38;5;221;48;5;180m▒\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;186m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;223m▒\033[38;5;136;48;5;144m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;224m░\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;144m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;137m▒\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;137m▓\033[38;5;94;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;223m░\033[38;5;178;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;186m▒\033[38;5;220;48;5;230m \033[38;5;220;48;5;230m \033[38;5;221;48;5;230m \033[38;5;94;48;5;186m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;214;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;187m▒\033[38;5;178;48;5;144m▓\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;224m░\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;172;48;5;95m▓\033[38;5;208;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;136;48;5;180m▒\033[38;5;220;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;172;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;180m▓\033[38;5;221;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;137m▓\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;187m▒\033[38;5;130;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;230m \033[38;5;136;48;5;187m▒\033[38;5;94;48;5;187m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;181m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;220;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;223m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;223m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;101m▒\033[38;5;221;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;181m▒\033[38;5;172;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;221;48;5;187m▒\033[38;5;221;48;5;187m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;130;48;5;180m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;221;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;178;48;5;186m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;94;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;130;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;253m▓\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;208;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;178;48;5;223m░\033[38;5;178;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;137m▒\033[38;5;221;48;5;101m▒\033[38;5;221;48;5;101m▒\033[38;5;221;48;5;137m▒\033[38;5;179;48;5;101m▒\033[38;5;130;48;5;144m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;224m░\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;208;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;137m▓\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;172;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;230m░\033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;186m░\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;94;48;5;101m▓\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;223m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;214;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;130;48;5;173m▒\033[38;5;224;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;144m▓\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;101m▓\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;186m░\033[38;5;136;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;178;48;5;223m▒\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;144m▓\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;179;48;5;187m▒\033[38;5;214;48;5;137m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;179m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;214;48;5;173m▒\033[38;5;221;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;220;48;5;181m▓\033[38;5;178;48;5;223m▒\033[38;5;94;48;5;101m▓\033[38;5;94;48;5;137m▓\033[38;5;214;48;5;144m▒\033[38;5;214;48;5;144m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;178;48;5;186m▒\033[38;5;220;48;5;180m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;187m▒\033[38;5;178;48;5;101m▓\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;143m▓\033[38;5;178;48;5;180m▒\033[38;5;94;48;5;144m▓\033[38;5;214;48;5;144m▓\033[38;5;221;48;5;144m▓\033[38;5;94;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;230m \033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;143m▒\033[38;5;221;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;137m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;214;48;5;223m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;224m▒\033[38;5;178;48;5;144m▓\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;186m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;255m▒\033[38;5;214;48;5;249m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;221;48;5;224m▒\033[38;5;221;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;187;48;5;187m▒\033[38;5;220;48;5;187m▓\033[38;5;179;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;214;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;230m░\033[38;5;179;48;5;144m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;255m░\033[38;5;136;48;5;187m▓\033[38;5;178;48;5;253m▒\033[38;5;230;48;5;230m \033[38;5;94;48;5;187m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;187m▒\033[38;5;179;48;5;187m▒\033[38;5;179;48;5;187m▒\033[38;5;94;48;5;230m░\033[38;5;230;48;5;231m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;254m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;223m░\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;223m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;179m▒\033[38;5;214;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;180m░\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;187m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;94;48;5;143m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;186m░\033[38;5;94;48;5;180m▒\033[38;5;136;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;224m▒\033[38;5;221;48;5;144m▓\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;220;48;5;180m▒\033[38;5;220;48;5;179m▒\033[38;5;220;48;5;143m▒\033[38;5;222;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;187m▒\033[38;5;179;48;5;179m▒\033[38;5;221;48;5;179m▒\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;214;48;5;180m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;144m▓\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;144m▒\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;179;48;5;186m▒\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;187m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;172;48;5;187m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;230m \033[38;5;172;48;5;180m▒\033[38;5;94;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;223m░\033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;187m▒\033[38;5;179;48;5;144m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;220;48;5;187m▒\033[38;5;185;48;5;229m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;187m▒\033[38;5;136;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;144m▓\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;221;48;5;230m \033[38;5;220;48;5;230m▒\033[38;5;186;48;5;230m▒\033[38;5;148;48;5;230m▒\033[38;5;148;48;5;255m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");

				$display("\n\033[1;32mCongratulations! Your critical path is below 3.5!\033[m\n");
			end
			else begin
				$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;223m▒\033[38;5;220;48;5;144m▓\033[38;5;178;48;5;137m▓\033[38;5;178;48;5;143m▓\033[38;5;178;48;5;180m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;94;48;5;186m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;180;48;5;180m▒\033[38;5;180;48;5;180m▒\033[38;5;208;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;186m░\033[38;5;172;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;221;48;5;229m \033[38;5;220;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;130;48;5;222m░\033[38;5;215;48;5;216m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;179m▒\033[38;5;208;48;5;179m▒\033[38;5;208;48;5;179m▒\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;130;48;5;179m▒\033[38;5;180;48;5;180m▒\033[38;5;202;48;5;181m▒\033[38;5;130;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;221;48;5;223m \033[38;5;130;48;5;216m░\033[38;5;166;48;5;216m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;179m▒\033[38;5;166;48;5;179m▒\033[38;5;180;48;5;179m▒\033[38;5;208;48;5;179m▒\033[38;5;166;48;5;179m▒\033[38;5;180;48;5;179m▒\033[38;5;180;48;5;137m▒\033[38;5;137;48;5;137m▓\033[38;5;130;48;5;187m▒\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;230m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;179m░\033[38;5;215;48;5;179m░\033[38;5;166;48;5;179m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;187m▒\033[38;5;222;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;221;48;5;229m \033[38;5;172;48;5;223m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;221m \033[38;5;130;48;5;215m░\033[38;5;180;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;215;48;5;179m░\033[38;5;208;48;5;179m░\033[38;5;215;48;5;179m░\033[38;5;180;48;5;179m░\033[38;5;180;48;5;179m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;185;48;5;230m░\033[38;5;220;48;5;187m▒\033[38;5;172;48;5;223m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;180;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;216m░\033[38;5;166;48;5;216m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;180m▒\033[38;5;166;48;5;224m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;187;48;5;187m▓\033[38;5;220;48;5;144m▓\033[38;5;130;48;5;222m \033[38;5;130;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;202;48;5;215m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;130m▒\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;136;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;187;48;5;253m▒\033[38;5;190;48;5;101m▓\033[38;5;143;48;5;240m▒\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;222m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;215;48;5;215m \033[38;5;215;48;5;215m \033[38;5;215;48;5;216m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;166;48;5;179m░\033[38;5;166;48;5;216m░\033[38;5;202;48;5;216m \033[38;5;202;48;5;215m \033[38;5;202;48;5;215m \033[38;5;202;48;5;209m \033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;130m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;130m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;137m▒\033[38;5;130;48;5;179m▒\033[38;5;221;48;5;229m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;144;48;5;252m▓\033[38;5;101;48;5;102m▓\033[38;5;178;48;5;245m▓\033[38;5;166;48;5;180m░\033[38;5;166;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;137m▒\033[38;5;76;48;5;244m▓\033[38;5;74;48;5;66m▓\033[38;5;67;48;5;238m▓\033[38;5;209;48;5;237m▓\033[38;5;166;48;5;237m▓\033[38;5;202;48;5;237m▒\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m \033[38;5;202;48;5;215m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;130m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;180m▒\033[38;5;220;48;5;230m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;180;48;5;181m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;209;48;5;131m▒\033[38;5;209;48;5;131m▒\033[38;5;204;48;5;138m▓\033[38;5;146;48;5;140m▒\033[38;5;68;48;5;110m▒\033[38;5;26;48;5;110m▒\033[38;5;67;48;5;247m▓\033[38;5;247;48;5;247m▓\033[38;5;202;48;5;144m▓\033[38;5;130;48;5;216m░\033[38;5;172;48;5;222m \033[38;5;222;48;5;222m \033[38;5;94;48;5;222m \033[38;5;221;48;5;222m \033[38;5;94;48;5;222m \033[38;5;222;48;5;222m \033[38;5;130;48;5;216m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;167m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;94;48;5;186m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;223;48;5;224m \033[38;5;137;48;5;138m▒\033[38;5;208;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;173m▒\033[38;5;130;48;5;180m▒\033[38;5;144;48;5;249m▓\033[38;5;66;48;5;7m▓\033[38;5;130;48;5;252m▓\033[38;5;172;48;5;223m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;222;48;5;222m \033[38;5;94;48;5;222m \033[38;5;178;48;5;222m \033[38;5;220;48;5;228m \033[38;5;220;48;5;229m \033[38;5;220;48;5;228m \033[38;5;221;48;5;222m \033[38;5;222;48;5;221m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;178;48;5;186m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;179;48;5;181m▓\033[38;5;172;48;5;138m▓\033[38;5;172;48;5;101m▓\033[38;5;130;48;5;95m▒\033[38;5;137;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;215;48;5;215m░\033[38;5;130;48;5;216m░\033[38;5;178;48;5;187m▒\033[38;5;25;48;5;251m▓\033[38;5;45;48;5;251m▓\033[38;5;190;48;5;187m▒\033[38;5;178;48;5;223m░\033[38;5;94;48;5;223m \033[38;5;94;48;5;223m░\033[38;5;221;48;5;223m░\033[38;5;178;48;5;229m \033[38;5;220;48;5;229m \033[38;5;220;48;5;229m \033[38;5;220;48;5;229m \033[38;5;136;48;5;229m \033[38;5;94;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;137m▓\033[38;5;166;48;5;144m▓\033[38;5;202;48;5;224m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;187m▓\033[38;5;220;48;5;245m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;136;48;5;95m▓\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;101m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;173m▒\033[38;5;130;48;5;179m░\033[38;5;208;48;5;215m░\033[38;5;208;48;5;216m░\033[38;5;130;48;5;216m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;216m░\033[38;5;214;48;5;186m▒\033[38;5;74;48;5;152m▓\033[38;5;33;48;5;110m▒\033[38;5;35;48;5;152m▒\033[38;5;149;48;5;187m▒\033[38;5;190;48;5;187m▒\033[38;5;220;48;5;224m▒\033[38;5;136;48;5;230m░\033[38;5;221;48;5;230m░\033[38;5;172;48;5;230m \033[38;5;172;48;5;230m \033[38;5;94;48;5;230m \033[38;5;221;48;5;230m \033[38;5;221;48;5;223m \033[38;5;214;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;173;48;5;180m▒\033[38;5;130;48;5;224m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;144;48;5;231m▓\033[38;5;101;48;5;247m▓\033[38;5;101;48;5;239m▓\033[38;5;143;48;5;239m▓\033[38;5;143;48;5;238m▒\033[38;5;186;48;5;58m▒\033[38;5;220;48;5;239m▒\033[38;5;221;48;5;95m▓\033[38;5;94;48;5;101m▓\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m░\033[38;5;130;48;5;179m░\033[38;5;130;48;5;179m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;70;48;5;249m▓\033[38;5;32;48;5;109m▓\033[38;5;72;48;5;250m▓\033[38;5;148;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;130;48;5;223m░\033[38;5;172;48;5;224m░\033[38;5;172;48;5;224m \033[38;5;222;48;5;230m \033[38;5;214;48;5;230m \033[38;5;222;48;5;224m \033[38;5;94;48;5;223m \033[38;5;221;48;5;223m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;209;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;172;48;5;180m▒\033[38;5;221;48;5;230m░\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;101;48;5;248m▓\033[38;5;220;48;5;239m▓\033[38;5;101;48;5;238m▓\033[38;5;143;48;5;236m▒\033[38;5;185;48;5;236m▒\033[38;5;58;48;5;58m░\033[38;5;58;48;5;58m░\033[38;5;178;48;5;58m▒\033[38;5;179;48;5;95m▓\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;220;48;5;101m▓\033[38;5;144;48;5;101m▓\033[38;5;136;48;5;137m▓\033[38;5;94;48;5;144m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;223m░\033[38;5;94;48;5;223m░\033[38;5;214;48;5;223m░\033[38;5;214;48;5;223m░\033[38;5;172;48;5;223m \033[38;5;222;48;5;223m \033[38;5;214;48;5;223m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;216m \033[38;5;130;48;5;216m \033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;187m▒\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;190;48;5;188m▓\033[38;5;148;48;5;240m▓\033[38;5;143;48;5;235m▓\033[38;5;143;48;5;236m▒\033[38;5;186;48;5;236m▒\033[38;5;186;48;5;236m▒\033[38;5;178;48;5;237m▒\033[38;5;221;48;5;240m▓\033[38;5;94;48;5;101m▓\033[38;5;179;48;5;144m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;137m▒\033[38;5;221;48;5;101m▒\033[38;5;136;48;5;58m░\033[38;5;221;48;5;58m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;223m░\033[38;5;94;48;5;223m \033[38;5;136;48;5;223m \033[38;5;221;48;5;223m \033[38;5;94;48;5;223m \033[38;5;94;48;5;223m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;208;48;5;173m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;185;48;5;230m░\033[38;5;101;48;5;249m▓\033[38;5;101;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;144m▓\033[38;5;179;48;5;144m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;94m▒\033[38;5;136;48;5;94m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;214;48;5;223m░\033[38;5;221;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;216m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;106;48;5;255m▒\033[38;5;190;48;5;188m▓\033[38;5;101;48;5;7m▓\033[38;5;220;48;5;249m▓\033[38;5;178;48;5;249m▓\033[38;5;178;48;5;144m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;137m▓\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;223m░\033[38;5;214;48;5;223m \033[38;5;94;48;5;223m \033[38;5;94;48;5;223m \033[38;5;94;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;223m \033[38;5;94;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;222m \033[38;5;130;48;5;216m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;208;48;5;173m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;186m▒\033[38;5;229;48;5;229m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;187;48;5;187m▒\033[38;5;220;48;5;144m▓\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;222;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;214;48;5;223m \033[38;5;214;48;5;223m \033[38;5;94;48;5;223m \033[38;5;94;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;222m \033[38;5;214;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;222m \033[38;5;130;48;5;216m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;214;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;190;48;5;230m░\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;214;48;5;223m░\033[38;5;214;48;5;223m░\033[38;5;94;48;5;223m \033[38;5;94;48;5;223m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;222m \033[38;5;208;48;5;216m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;202;48;5;215m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;209;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;223;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;64;48;5;230m \033[38;5;220;48;5;187m▒\033[38;5;94;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;214;48;5;223m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;130;48;5;222m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;173m░\033[38;5;209;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;179m▒\033[38;5;180;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;154;48;5;230m░\033[38;5;136;48;5;187m▒\033[38;5;172;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;223;48;5;223m \033[38;5;223;48;5;223m░\033[38;5;208;48;5;223m░\033[38;5;208;48;5;223m░\033[38;5;208;48;5;223m \033[38;5;130;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;221m░\033[38;5;172;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;173m▒\033[38;5;208;48;5;179m▒\033[38;5;172;48;5;223m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m░\033[38;5;172;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;130;48;5;223m \033[38;5;208;48;5;223m \033[38;5;223;48;5;223m░\033[38;5;223;48;5;223m░\033[38;5;223;48;5;223m░\033[38;5;223;48;5;223m░\033[38;5;223;48;5;223m░\033[38;5;208;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;214;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;222;48;5;221m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;208;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;209;48;5;173m░\033[38;5;209;48;5;173m░\033[38;5;209;48;5;173m░\033[38;5;209;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;130;48;5;180m▒\033[38;5;214;48;5;223m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;230m \033[38;5;208;48;5;224m░\033[38;5;130;48;5;144m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;137;48;5;235m▓\033[38;5;137;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;172;48;5;235m▓\033[38;5;172;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;172;48;5;234m▒\033[38;5;172;48;5;95m▒\033[38;5;130;48;5;179m░\033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;131m▒\033[38;5;202;48;5;233m░\033[38;5;202;48;5;233m░\033[38;5;202;48;5;233m \033[38;5;216;48;5;233m \033[38;5;216;48;5;233m \033[38;5;202;48;5;235m░\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;209m \033[38;5;202;48;5;209m \033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m \033[38;5;202;48;5;173m▒\033[38;5;202;48;5;238m▒\033[38;5;202;48;5;234m░\033[38;5;202;48;5;234m░\033[38;5;202;48;5;234m░\033[38;5;166;48;5;234m░\033[38;5;166;48;5;238m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;237m▒\033[38;5;166;48;5;233m░\033[38;5;215;48;5;233m░\033[38;5;166;48;5;233m░\033[38;5;166;48;5;233m░\033[38;5;166;48;5;238m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;172;48;5;180m▒\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;215m░\033[38;5;202;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;208;48;5;179m▒\033[38;5;172;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;246;48;5;246m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;242m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;130;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;239m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;130;48;5;180m▒\033[38;5;220;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;130;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;243;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;179;48;5;233m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;239m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;94m▒\033[38;5;202;48;5;130m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;180m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;243;48;5;242m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;239m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;94m▒\033[38;5;173;48;5;94m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;250;48;5;250m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;239;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;239m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;94m▒\033[38;5;173;48;5;94m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;95m▒\033[38;5;172;48;5;101m▓\033[38;5;94;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;179;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;241;48;5;241m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;239m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;130m▒\033[38;5;173;48;5;130m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;95m▒\033[38;5;137;48;5;95m▓\033[38;5;130;48;5;138m▓\033[38;5;202;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;253;48;5;253m▓\033[38;5;254;48;5;254m▓\033[38;5;253;48;5;253m▓\033[38;5;253;48;5;253m▓\033[38;5;253;48;5;253m▓\033[38;5;254;48;5;254m▓\033[38;5;253;48;5;253m▓\033[38;5;236;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;233;48;5;233m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;235m▒\033[38;5;166;48;5;58m▒\033[38;5;202;48;5;58m▒\033[38;5;202;48;5;58m▒\033[38;5;202;48;5;58m▒\033[38;5;202;48;5;95m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;137;48;5;95m▓\033[38;5;208;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;101;48;5;242m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;252;48;5;251m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;241;48;5;241m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;232m \033[38;5;202;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;130;48;5;101m▓\033[38;5;222;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;242m▓\033[38;5;179;48;5;245m▓\033[38;5;179;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;246;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;236;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;243;48;5;243m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;236;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;246;48;5;246m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;239m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;172;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;172;48;5;242m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;235;48;5;235m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;237m▓\033[38;5;214;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;250;48;5;250m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;252m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;239m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;208;48;5;173m▒\033[38;5;179;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;250m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;234m▓\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;223m░\033[38;5;214;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;179;48;5;95m▓\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;179;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;95m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;179;48;5;144m▓\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;94;48;5;187m▒\033[38;5;94;48;5;101m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;235m▓\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;186m▒\033[38;5;94;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;95m▓\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;220;48;5;232m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;233m▒\033[38;5;208;48;5;237m▒\033[38;5;180;48;5;232m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;130;48;5;233m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;214;48;5;137m▓\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;223m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;221m░\033[38;5;222;48;5;215m░\033[38;5;179;48;5;215m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;216m \033[38;5;130;48;5;216m \033[38;5;208;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;208;48;5;179m░\033[38;5;180;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;214;48;5;144m▓\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;223m░\033[38;5;214;48;5;186m░\033[38;5;222;48;5;221m░\033[38;5;172;48;5;221m░\033[38;5;172;48;5;221m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;179;48;5;180m░\033[38;5;179;48;5;180m░\033[38;5;179;48;5;180m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;172;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;186m░\033[38;5;179;48;5;216m░\033[38;5;172;48;5;221m \033[38;5;172;48;5;221m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;180;48;5;179m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▓\033[38;5;130;48;5;137m▓\033[38;5;222;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;186m▒\033[38;5;179;48;5;215m░\033[38;5;172;48;5;221m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;130;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;137;48;5;131m▒\033[38;5;208;48;5;101m▓\033[38;5;208;48;5;138m▓\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;186m▒\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;137;48;5;137m▓\033[38;5;137;48;5;137m▓\033[38;5;209;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;186m▒\033[38;5;222;48;5;222m░\033[38;5;214;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;95m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;130;48;5;137m▓\033[38;5;130;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;222;48;5;222m \033[38;5;94;48;5;222m \033[38;5;222;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;216m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;179m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;180m▒\033[38;5;208;48;5;224m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;216m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;202;48;5;131m▒\033[38;5;180;48;5;95m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;137;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;180m▒\033[38;5;221;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;229;48;5;229m \033[38;5;94;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m░\033[38;5;214;48;5;180m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;94m▒\033[38;5;179;48;5;94m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;130;48;5;94m▒\033[38;5;179;48;5;58m░\033[38;5;179;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;130;48;5;95m▒\033[38;5;130;48;5;95m▒\033[38;5;130;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;137;48;5;137m▒\033[38;5;137;48;5;137m▓\033[38;5;130;48;5;180m▒\033[38;5;136;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;172;48;5;221m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;101m▒\033[38;5;221;48;5;101m▒\033[38;5;221;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;208;48;5;95m▒\033[38;5;172;48;5;58m░\033[38;5;179;48;5;58m░\033[38;5;179;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;208;48;5;95m▒\033[38;5;130;48;5;95m▒\033[38;5;208;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;208;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;137m▓\033[38;5;130;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;220;48;5;230m \033[38;5;220;48;5;223m░\033[38;5;220;48;5;187m▒\033[38;5;186;48;5;187m▒\033[38;5;186;48;5;186m▒\033[38;5;186;48;5;186m▒\033[38;5;186;48;5;186m▒\033[38;5;186;48;5;186m▒\033[38;5;186;48;5;186m▒\033[38;5;220;48;5;185m▒\033[38;5;94;48;5;221m░\033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;186m▒\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;137m▒\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;101m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;137m▓\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;221m \033[38;5;172;48;5;221m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;180;48;5;95m▒\033[38;5;130;48;5;58m▒\033[38;5;179;48;5;58m░\033[38;5;94;48;5;58m▒\033[38;5;214;48;5;58m▒\033[38;5;179;48;5;58m▒\033[38;5;214;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;180m▒\033[38;5;136;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;136;48;5;230m░\033[38;5;136;48;5;224m▒\033[38;5;220;48;5;223m▒\033[38;5;220;48;5;223m▒\033[38;5;220;48;5;223m░\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;186;48;5;186m▒\033[38;5;220;48;5;180m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;94m▒\033[38;5;221;48;5;58m░\033[38;5;179;48;5;95m▒\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;221m \033[38;5;130;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;208;48;5;95m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;58m░\033[38;5;179;48;5;58m▒\033[38;5;179;48;5;58m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;94;48;5;95m▒\033[38;5;94;48;5;95m▓\033[38;5;214;48;5;144m▓\033[38;5;136;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;136;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;185;48;5;223m░\033[38;5;185;48;5;223m▒\033[38;5;185;48;5;187m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;178;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;220;48;5;144m▒\033[38;5;178;48;5;144m▓\033[38;5;178;48;5;144m▓\033[38;5;178;48;5;186m▒\033[38;5;94;48;5;223m░\033[38;5;221;48;5;229m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;95m▒\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;238m▒\033[38;5;179;48;5;240m▓\033[38;5;172;48;5;144m▓\033[38;5;220;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;144;48;5;253m▓\033[38;5;220;48;5;101m▓\033[38;5;187;48;5;150m▓\033[38;5;186;48;5;187m▒\033[38;5;143;48;5;144m▒\033[38;5;143;48;5;101m▓\033[38;5;144;48;5;143m▓\033[38;5;143;48;5;144m▓\033[38;5;187;48;5;180m▓\033[38;5;187;48;5;187m▒\033[38;5;185;48;5;193m▒\033[38;5;230;48;5;230m░\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;130;48;5;223m \033[38;5;130;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;222;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;95m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;239m▒\033[38;5;172;48;5;239m▒\033[38;5;179;48;5;239m▒\033[38;5;179;48;5;240m▒\033[38;5;172;48;5;95m▓\033[38;5;172;48;5;137m▓\033[38;5;172;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;185;48;5;230m▒\033[38;5;187;48;5;254m▓\033[38;5;185;48;5;230m░\033[38;5;187;48;5;253m▓\033[38;5;144;48;5;187m▓\033[38;5;144;48;5;187m▓\033[38;5;186;48;5;255m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;220;48;5;229m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m░\033[38;5;172;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;172;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;131m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;238m▒\033[38;5;172;48;5;239m▒\033[38;5;172;48;5;239m▓\033[38;5;172;48;5;95m▓\033[38;5;172;48;5;101m▓\033[38;5;130;48;5;144m▓\033[38;5;223;48;5;224m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;220;48;5;229m \033[38;5;172;48;5;180m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;222;48;5;222m \033[38;5;214;48;5;221m \033[38;5;214;48;5;221m \033[38;5;172;48;5;221m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;178;48;5;137m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;94;48;5;223m░\033[38;5;179;48;5;223m░\033[38;5;179;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;179;48;5;223m░\033[38;5;94;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;94m▒\033[38;5;179;48;5;58m░\033[38;5;94;48;5;58m▒\033[38;5;221;48;5;58m▒\033[38;5;179;48;5;237m▒\033[38;5;172;48;5;95m▓\033[38;5;172;48;5;181m▓\033[38;5;220;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;230m \033[38;5;178;48;5;223m░\033[38;5;221;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;214;48;5;221m \033[38;5;214;48;5;221m░\033[38;5;222;48;5;221m░\033[38;5;222;48;5;221m░\033[38;5;172;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;223m░\033[38;5;94;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;179;48;5;223m░\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;130;48;5;101m▓\033[38;5;179;48;5;187m▒\033[38;5;220;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;136;48;5;229m░\033[38;5;221;48;5;223m░\033[38;5;136;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;222;48;5;221m░\033[38;5;222;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;186m░\033[38;5;172;48;5;223m░\033[38;5;130;48;5;181m▒\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;181m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;223m░\033[38;5;222;48;5;224m \033[38;5;214;48;5;223m░\033[38;5;222;48;5;230m \033[38;5;222;48;5;230m \033[38;5;172;48;5;224m \033[38;5;172;48;5;224m \033[38;5;222;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;179;48;5;223m░\033[38;5;94;48;5;223m▒\033[38;5;221;48;5;187m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;144m▒\033[38;5;221;48;5;143m▒\033[38;5;172;48;5;180m▒\033[38;5;130;48;5;216m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▓\033[38;5;137;48;5;137m▓\033[38;5;166;48;5;144m▓\033[38;5;166;48;5;188m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;223m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;178;48;5;230m \033[38;5;179;48;5;186m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;216m░\033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;137;48;5;137m▓\033[38;5;208;48;5;138m▓\033[38;5;178;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;231m \033[38;5;220;48;5;144m▓\033[38;5;220;48;5;101m▓\033[38;5;178;48;5;137m▓\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;179;48;5;180m░\033[38;5;179;48;5;180m░\033[38;5;222;48;5;222m░\033[38;5;94;48;5;222m \033[38;5;136;48;5;222m \033[38;5;136;48;5;222m \033[38;5;178;48;5;222m \033[38;5;178;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;220;48;5;222m░\033[38;5;220;48;5;222m░\033[38;5;220;48;5;186m░\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;222;48;5;223m \033[38;5;130;48;5;222m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;180m▓\033[38;5;172;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;231m \033[38;5;94;48;5;187m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m \033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;221;48;5;222m \033[38;5;136;48;5;222m \033[38;5;178;48;5;222m \033[38;5;178;48;5;222m \033[38;5;178;48;5;222m \033[38;5;220;48;5;222m░\033[38;5;220;48;5;228m░\033[38;5;185;48;5;186m░\033[38;5;229;48;5;229m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;223m \033[38;5;130;48;5;222m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;214;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;230m \033[38;5;94;48;5;187m▒\033[38;5;221;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;221;48;5;222m \033[38;5;221;48;5;222m \033[38;5;221;48;5;222m \033[38;5;136;48;5;222m \033[38;5;136;48;5;222m \033[38;5;178;48;5;222m░\033[38;5;220;48;5;222m░\033[38;5;229;48;5;229m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;178;48;5;229m \033[38;5;172;48;5;222m \033[38;5;172;48;5;221m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;230m \033[38;5;178;48;5;223m░\033[38;5;136;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;222m \033[38;5;221;48;5;222m \033[38;5;221;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;222;48;5;222m \033[38;5;221;48;5;223m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;172;48;5;223m \033[38;5;130;48;5;222m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;221;48;5;224m░\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;94;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;172;48;5;223m \033[38;5;130;48;5;216m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;172;48;5;222m \033[38;5;130;48;5;216m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;220;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;229m \033[38;5;130;48;5;222m \033[38;5;130;48;5;216m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;181m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;94;48;5;223m \033[38;5;172;48;5;222m \033[38;5;130;48;5;216m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;180;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;94;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;94;48;5;223m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;180;48;5;179m▒\033[38;5;166;48;5;216m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;214;48;5;223m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;208;48;5;179m░\033[38;5;180;48;5;179m▒\033[38;5;166;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m░\033[38;5;94;48;5;187m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;222m░\033[38;5;130;48;5;222m░\033[38;5;130;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;215m \033[38;5;166;48;5;215m \033[38;5;215;48;5;179m░\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;172;48;5;224m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;181m▓\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;216m░\033[38;5;172;48;5;180m░\033[38;5;130;48;5;179m░\033[38;5;130;48;5;179m░\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;180m▒\033[38;5;94;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;144m▓\033[38;5;172;48;5;101m▓\033[38;5;172;48;5;144m▓\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;143m▓\033[38;5;178;48;5;95m▓\033[38;5;220;48;5;137m▓\033[38;5;220;48;5;223m▒\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
			end

			if(err3 == 0) begin

			end
			else if(err4 == 0)
				$display("\n\033[1;32mCongratulations! Your critical path is below 4!\033[m\n");
			else if(err5 == 0)
				$display("\n\033[1;32mCongratulations! Your critical path is below 4.5!\033[m\n");
			else if(err6 == 0)
				$display("\n\033[1;32mCongratulations! Your critical path is below 5!\033[m\n");
			else if(err7 == 0)
				$display("\n\033[1;32mCongratulations! Your critical path is below 5.5!\033[m\n");
			else if(err10 == 0)
				$display("\n\033[1;32mCongratulations! Your critical path is below 6!\033[m\n");
			else if(err20 == 0)
				$display("\n\033[1;32mCongratulations! Your score is 40!\033[m\n");
			else begin
			   $display("\nThere are %d errors.\n", err20);
			   $display("Your score is %g.\n", 40-err20/25);
			end


			$finish;
		end
		if (err20>100)begin
			$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;223m▒\033[38;5;220;48;5;144m▓\033[38;5;178;48;5;137m▓\033[38;5;178;48;5;143m▓\033[38;5;178;48;5;180m▒\033[38;5;178;48;5;187m▒\033[38;5;220;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;94;48;5;186m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;180;48;5;180m▒\033[38;5;180;48;5;180m▒\033[38;5;208;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;186m░\033[38;5;172;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;221;48;5;229m \033[38;5;220;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;130;48;5;222m░\033[38;5;215;48;5;216m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;179m▒\033[38;5;208;48;5;179m▒\033[38;5;208;48;5;179m▒\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;130;48;5;179m▒\033[38;5;180;48;5;180m▒\033[38;5;202;48;5;181m▒\033[38;5;130;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;221;48;5;223m \033[38;5;130;48;5;216m░\033[38;5;166;48;5;216m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;179m▒\033[38;5;166;48;5;179m▒\033[38;5;180;48;5;179m▒\033[38;5;208;48;5;179m▒\033[38;5;166;48;5;179m▒\033[38;5;180;48;5;179m▒\033[38;5;180;48;5;137m▒\033[38;5;137;48;5;137m▓\033[38;5;130;48;5;187m▒\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;230m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;179m░\033[38;5;215;48;5;179m░\033[38;5;166;48;5;179m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;187m▒\033[38;5;222;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;221;48;5;229m \033[38;5;172;48;5;223m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;221m \033[38;5;130;48;5;215m░\033[38;5;180;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;215;48;5;179m░\033[38;5;208;48;5;179m░\033[38;5;215;48;5;179m░\033[38;5;180;48;5;179m░\033[38;5;180;48;5;179m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;185;48;5;230m░\033[38;5;220;48;5;187m▒\033[38;5;172;48;5;223m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;180;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;216m░\033[38;5;166;48;5;216m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;180m▒\033[38;5;166;48;5;224m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;187;48;5;187m▓\033[38;5;220;48;5;144m▓\033[38;5;130;48;5;222m \033[38;5;130;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;202;48;5;215m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;130m▒\033[38;5;166;48;5;94m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;136;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;187;48;5;253m▒\033[38;5;190;48;5;101m▓\033[38;5;143;48;5;240m▒\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;222m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;215;48;5;215m \033[38;5;215;48;5;215m \033[38;5;215;48;5;216m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;166;48;5;179m░\033[38;5;166;48;5;216m░\033[38;5;202;48;5;216m \033[38;5;202;48;5;215m \033[38;5;202;48;5;215m \033[38;5;202;48;5;209m \033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;130m▒\033[38;5;202;48;5;94m▒\033[38;5;202;48;5;130m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;137m▒\033[38;5;130;48;5;179m▒\033[38;5;221;48;5;229m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;144;48;5;252m▓\033[38;5;101;48;5;102m▓\033[38;5;178;48;5;245m▓\033[38;5;166;48;5;180m░\033[38;5;166;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;137m▒\033[38;5;76;48;5;244m▓\033[38;5;74;48;5;66m▓\033[38;5;67;48;5;238m▓\033[38;5;209;48;5;237m▓\033[38;5;166;48;5;237m▓\033[38;5;202;48;5;237m▒\033[38;5;166;48;5;58m░\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m \033[38;5;202;48;5;215m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;130m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;180m▒\033[38;5;220;48;5;230m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;180;48;5;181m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;209;48;5;131m▒\033[38;5;209;48;5;131m▒\033[38;5;204;48;5;138m▓\033[38;5;146;48;5;140m▒\033[38;5;68;48;5;110m▒\033[38;5;26;48;5;110m▒\033[38;5;67;48;5;247m▓\033[38;5;247;48;5;247m▓\033[38;5;202;48;5;144m▓\033[38;5;130;48;5;216m░\033[38;5;172;48;5;222m \033[38;5;222;48;5;222m \033[38;5;94;48;5;222m \033[38;5;221;48;5;222m \033[38;5;94;48;5;222m \033[38;5;222;48;5;222m \033[38;5;130;48;5;216m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;167m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;94;48;5;186m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;223;48;5;224m \033[38;5;137;48;5;138m▒\033[38;5;208;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;173m▒\033[38;5;130;48;5;180m▒\033[38;5;144;48;5;249m▓\033[38;5;66;48;5;7m▓\033[38;5;130;48;5;252m▓\033[38;5;172;48;5;223m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;222;48;5;222m \033[38;5;94;48;5;222m \033[38;5;178;48;5;222m \033[38;5;220;48;5;228m \033[38;5;220;48;5;229m \033[38;5;220;48;5;228m \033[38;5;221;48;5;222m \033[38;5;222;48;5;221m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;178;48;5;186m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;179;48;5;181m▓\033[38;5;172;48;5;138m▓\033[38;5;172;48;5;101m▓\033[38;5;130;48;5;95m▒\033[38;5;137;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;215;48;5;215m░\033[38;5;130;48;5;216m░\033[38;5;178;48;5;187m▒\033[38;5;25;48;5;251m▓\033[38;5;45;48;5;251m▓\033[38;5;190;48;5;187m▒\033[38;5;178;48;5;223m░\033[38;5;94;48;5;223m \033[38;5;94;48;5;223m░\033[38;5;221;48;5;223m░\033[38;5;178;48;5;229m \033[38;5;220;48;5;229m \033[38;5;220;48;5;229m \033[38;5;220;48;5;229m \033[38;5;136;48;5;229m \033[38;5;94;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;137m▓\033[38;5;166;48;5;144m▓\033[38;5;202;48;5;224m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;187m▓\033[38;5;220;48;5;245m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;136;48;5;95m▓\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;101m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;173m▒\033[38;5;130;48;5;179m░\033[38;5;208;48;5;215m░\033[38;5;208;48;5;216m░\033[38;5;130;48;5;216m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;216m░\033[38;5;214;48;5;186m▒\033[38;5;74;48;5;152m▓\033[38;5;33;48;5;110m▒\033[38;5;35;48;5;152m▒\033[38;5;149;48;5;187m▒\033[38;5;190;48;5;187m▒\033[38;5;220;48;5;224m▒\033[38;5;136;48;5;230m░\033[38;5;221;48;5;230m░\033[38;5;172;48;5;230m \033[38;5;172;48;5;230m \033[38;5;94;48;5;230m \033[38;5;221;48;5;230m \033[38;5;221;48;5;223m \033[38;5;214;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;173;48;5;180m▒\033[38;5;130;48;5;224m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;144;48;5;231m▓\033[38;5;101;48;5;247m▓\033[38;5;101;48;5;239m▓\033[38;5;143;48;5;239m▓\033[38;5;143;48;5;238m▒\033[38;5;186;48;5;58m▒\033[38;5;220;48;5;239m▒\033[38;5;221;48;5;95m▓\033[38;5;94;48;5;101m▓\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m░\033[38;5;130;48;5;179m░\033[38;5;130;48;5;179m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;70;48;5;249m▓\033[38;5;32;48;5;109m▓\033[38;5;72;48;5;250m▓\033[38;5;148;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;130;48;5;223m░\033[38;5;172;48;5;224m░\033[38;5;172;48;5;224m \033[38;5;222;48;5;230m \033[38;5;214;48;5;230m \033[38;5;222;48;5;224m \033[38;5;94;48;5;223m \033[38;5;221;48;5;223m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;209;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;172;48;5;180m▒\033[38;5;221;48;5;230m░\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;101;48;5;248m▓\033[38;5;220;48;5;239m▓\033[38;5;101;48;5;238m▓\033[38;5;143;48;5;236m▒\033[38;5;185;48;5;236m▒\033[38;5;58;48;5;58m░\033[38;5;58;48;5;58m░\033[38;5;178;48;5;58m▒\033[38;5;179;48;5;95m▓\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;220;48;5;101m▓\033[38;5;144;48;5;101m▓\033[38;5;136;48;5;137m▓\033[38;5;94;48;5;144m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;223m░\033[38;5;94;48;5;223m░\033[38;5;214;48;5;223m░\033[38;5;214;48;5;223m░\033[38;5;172;48;5;223m \033[38;5;222;48;5;223m \033[38;5;214;48;5;223m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;216m \033[38;5;130;48;5;216m \033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;130;48;5;173m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;187m▒\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;190;48;5;188m▓\033[38;5;148;48;5;240m▓\033[38;5;143;48;5;235m▓\033[38;5;143;48;5;236m▒\033[38;5;186;48;5;236m▒\033[38;5;186;48;5;236m▒\033[38;5;178;48;5;237m▒\033[38;5;221;48;5;240m▓\033[38;5;94;48;5;101m▓\033[38;5;179;48;5;144m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;143m▒\033[38;5;214;48;5;137m▒\033[38;5;221;48;5;101m▒\033[38;5;136;48;5;58m░\033[38;5;221;48;5;58m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;143m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;214;48;5;223m░\033[38;5;94;48;5;223m \033[38;5;136;48;5;223m \033[38;5;221;48;5;223m \033[38;5;94;48;5;223m \033[38;5;94;48;5;223m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;208;48;5;173m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;185;48;5;230m░\033[38;5;101;48;5;249m▓\033[38;5;101;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;220;48;5;101m▓\033[38;5;136;48;5;101m▓\033[38;5;221;48;5;137m▓\033[38;5;94;48;5;144m▓\033[38;5;179;48;5;144m▒\033[38;5;179;48;5;143m▒\033[38;5;179;48;5;137m▒\033[38;5;214;48;5;137m▒\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;101m▒\033[38;5;94;48;5;94m▒\033[38;5;136;48;5;94m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;137m▓\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;214;48;5;223m░\033[38;5;221;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;216m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;106;48;5;255m▒\033[38;5;190;48;5;188m▓\033[38;5;101;48;5;7m▓\033[38;5;220;48;5;249m▓\033[38;5;178;48;5;249m▓\033[38;5;178;48;5;144m▓\033[38;5;136;48;5;101m▓\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;137m▓\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;137m▓\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;214;48;5;223m░\033[38;5;214;48;5;223m \033[38;5;94;48;5;223m \033[38;5;94;48;5;223m \033[38;5;94;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;223m \033[38;5;94;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;222m \033[38;5;130;48;5;216m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;208;48;5;173m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;94;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;186m▒\033[38;5;229;48;5;229m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;187;48;5;187m▒\033[38;5;220;48;5;144m▓\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;222;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;214;48;5;223m \033[38;5;214;48;5;223m \033[38;5;94;48;5;223m \033[38;5;94;48;5;223m \033[38;5;221;48;5;223m \033[38;5;221;48;5;222m \033[38;5;214;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;222m \033[38;5;130;48;5;216m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;214;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;190;48;5;230m░\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;214;48;5;223m░\033[38;5;214;48;5;223m░\033[38;5;94;48;5;223m \033[38;5;94;48;5;223m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;222m \033[38;5;208;48;5;216m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;202;48;5;215m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;209;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;223;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;64;48;5;230m \033[38;5;220;48;5;187m▒\033[38;5;94;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;214;48;5;223m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;130;48;5;222m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;173;48;5;167m▒\033[38;5;209;48;5;167m▒\033[38;5;209;48;5;173m░\033[38;5;209;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;179m▒\033[38;5;180;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;154;48;5;230m░\033[38;5;136;48;5;187m▒\033[38;5;172;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;223;48;5;223m \033[38;5;223;48;5;223m░\033[38;5;208;48;5;223m░\033[38;5;208;48;5;223m░\033[38;5;208;48;5;223m \033[38;5;130;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;221m░\033[38;5;172;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;209;48;5;167m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;173m▒\033[38;5;208;48;5;179m▒\033[38;5;172;48;5;223m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m░\033[38;5;172;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;130;48;5;223m \033[38;5;208;48;5;223m \033[38;5;223;48;5;223m░\033[38;5;223;48;5;223m░\033[38;5;223;48;5;223m░\033[38;5;223;48;5;223m░\033[38;5;223;48;5;223m░\033[38;5;208;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;214;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;222;48;5;221m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;208;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;209;48;5;173m░\033[38;5;209;48;5;173m░\033[38;5;209;48;5;173m░\033[38;5;209;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;216;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;130;48;5;180m▒\033[38;5;214;48;5;223m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;230m \033[38;5;208;48;5;224m░\033[38;5;130;48;5;144m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;137;48;5;235m▓\033[38;5;137;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;130;48;5;235m▓\033[38;5;172;48;5;235m▓\033[38;5;172;48;5;234m▒\033[38;5;179;48;5;234m▒\033[38;5;172;48;5;234m▒\033[38;5;172;48;5;95m▒\033[38;5;130;48;5;179m░\033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;131m▒\033[38;5;202;48;5;233m░\033[38;5;202;48;5;233m░\033[38;5;202;48;5;233m \033[38;5;216;48;5;233m \033[38;5;216;48;5;233m \033[38;5;202;48;5;235m░\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;209m \033[38;5;202;48;5;209m \033[38;5;202;48;5;209m░\033[38;5;202;48;5;209m \033[38;5;202;48;5;173m▒\033[38;5;202;48;5;238m▒\033[38;5;202;48;5;234m░\033[38;5;202;48;5;234m░\033[38;5;202;48;5;234m░\033[38;5;166;48;5;234m░\033[38;5;166;48;5;238m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;237m▒\033[38;5;166;48;5;233m░\033[38;5;215;48;5;233m░\033[38;5;166;48;5;233m░\033[38;5;166;48;5;233m░\033[38;5;166;48;5;238m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;172;48;5;180m▒\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;215m░\033[38;5;202;48;5;16m \033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;208;48;5;179m▒\033[38;5;172;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;244m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;246;48;5;246m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;242;48;5;242m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;130;48;5;95m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;239m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;130;48;5;180m▒\033[38;5;220;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;130;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;243;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;179;48;5;233m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;239m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;94m▒\033[38;5;202;48;5;130m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;180m▒\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;243;48;5;242m▓\033[38;5;188;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;248;48;5;248m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;239m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;94m▒\033[38;5;173;48;5;94m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;250;48;5;250m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;239;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;239m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;94m▒\033[38;5;173;48;5;94m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;95m▒\033[38;5;172;48;5;101m▓\033[38;5;94;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;179;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;238;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;237;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;233;48;5;233m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;241;48;5;241m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;239m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;130m▒\033[38;5;173;48;5;130m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;95m▒\033[38;5;137;48;5;95m▓\033[38;5;130;48;5;138m▓\033[38;5;202;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;253;48;5;253m▓\033[38;5;254;48;5;254m▓\033[38;5;253;48;5;253m▓\033[38;5;253;48;5;253m▓\033[38;5;253;48;5;253m▓\033[38;5;254;48;5;254m▓\033[38;5;253;48;5;253m▓\033[38;5;236;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;233;48;5;233m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;254;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;253;48;5;188m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;235m▒\033[38;5;166;48;5;58m▒\033[38;5;202;48;5;58m▒\033[38;5;202;48;5;58m▒\033[38;5;202;48;5;58m▒\033[38;5;202;48;5;95m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;137;48;5;95m▓\033[38;5;208;48;5;145m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;101;48;5;242m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;252;48;5;251m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;241;48;5;241m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;232m \033[38;5;202;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;130m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;130;48;5;101m▓\033[38;5;222;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;243m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;242m▓\033[38;5;179;48;5;245m▓\033[38;5;179;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;246;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;236;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;243;48;5;243m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;236;48;5;236m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;251;48;5;251m▓\033[38;5;246;48;5;246m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;166;48;5;239m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;172;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;172;48;5;242m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;247;48;5;247m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;234m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;235;48;5;235m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;240;48;5;240m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;214;48;5;237m▓\033[38;5;214;48;5;235m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;250;48;5;250m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;254;48;5;254m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;253;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;188;48;5;252m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;239m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;208;48;5;173m▒\033[38;5;179;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;250m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;234m▓\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;223m░\033[38;5;214;48;5;237m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;179;48;5;95m▓\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;179;48;5;234m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;202;48;5;95m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;179;48;5;144m▓\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;94;48;5;187m▒\033[38;5;94;48;5;101m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;235m▓\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;186m▒\033[38;5;94;48;5;239m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;94;48;5;95m▓\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;238m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;220;48;5;232m▒\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;172;48;5;233m▒\033[38;5;208;48;5;237m▒\033[38;5;180;48;5;232m░\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;16;48;5;16m▓\033[38;5;130;48;5;233m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;214;48;5;137m▓\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;223m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;221m░\033[38;5;222;48;5;215m░\033[38;5;179;48;5;215m░\033[38;5;179;48;5;179m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;216m \033[38;5;130;48;5;216m \033[38;5;208;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;208;48;5;179m░\033[38;5;180;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;173;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;214;48;5;144m▓\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;223m░\033[38;5;214;48;5;186m░\033[38;5;222;48;5;221m░\033[38;5;172;48;5;221m░\033[38;5;172;48;5;221m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;179;48;5;180m░\033[38;5;179;48;5;180m░\033[38;5;179;48;5;180m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;179;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;172;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;186m░\033[38;5;179;48;5;216m░\033[38;5;172;48;5;221m \033[38;5;172;48;5;221m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;180;48;5;179m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;202;48;5;131m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▓\033[38;5;130;48;5;137m▓\033[38;5;222;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;186m▒\033[38;5;179;48;5;215m░\033[38;5;172;48;5;221m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;130;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;137;48;5;131m▒\033[38;5;208;48;5;101m▓\033[38;5;208;48;5;138m▓\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;186m▒\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;94m▒\033[38;5;166;48;5;95m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;137;48;5;137m▓\033[38;5;137;48;5;137m▓\033[38;5;209;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;186m▒\033[38;5;222;48;5;222m░\033[38;5;214;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;180m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;216m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;166;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;95m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;130;48;5;137m▓\033[38;5;130;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;222;48;5;222m \033[38;5;94;48;5;222m \033[38;5;222;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;216m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;179m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;131m▒\033[38;5;166;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;130;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;166;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;180m▒\033[38;5;208;48;5;224m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;221;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;222;48;5;222m \033[38;5;172;48;5;216m░\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;179;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;173;48;5;173m▒\033[38;5;202;48;5;131m▒\033[38;5;180;48;5;95m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m░\033[38;5;208;48;5;58m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;94m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;137;48;5;137m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;180m▒\033[38;5;221;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;229;48;5;229m \033[38;5;94;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m░\033[38;5;214;48;5;180m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;137m▒\033[38;5;94;48;5;101m▒\033[38;5;214;48;5;94m▒\033[38;5;179;48;5;94m▒\033[38;5;179;48;5;95m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;173;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;137m▒\033[38;5;180;48;5;131m▒\033[38;5;130;48;5;94m▒\033[38;5;179;48;5;58m░\033[38;5;179;48;5;58m░\033[38;5;172;48;5;58m░\033[38;5;130;48;5;58m▒\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;130;48;5;95m▒\033[38;5;130;48;5;95m▒\033[38;5;130;48;5;95m▒\033[38;5;180;48;5;95m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;166;48;5;131m▒\033[38;5;137;48;5;137m▒\033[38;5;137;48;5;137m▓\033[38;5;130;48;5;180m▒\033[38;5;136;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;220;48;5;230m░\033[38;5;220;48;5;187m▒\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;172;48;5;221m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;101m▒\033[38;5;221;48;5;101m▒\033[38;5;221;48;5;101m▒\033[38;5;179;48;5;101m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;202;48;5;209m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m░\033[38;5;202;48;5;173m▒\033[38;5;202;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;208;48;5;95m▒\033[38;5;172;48;5;58m░\033[38;5;179;48;5;58m░\033[38;5;179;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;208;48;5;95m▒\033[38;5;130;48;5;95m▒\033[38;5;208;48;5;131m▒\033[38;5;180;48;5;131m▒\033[38;5;208;48;5;131m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;137m▓\033[38;5;130;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;220;48;5;230m \033[38;5;220;48;5;223m░\033[38;5;220;48;5;187m▒\033[38;5;186;48;5;187m▒\033[38;5;186;48;5;186m▒\033[38;5;186;48;5;186m▒\033[38;5;186;48;5;186m▒\033[38;5;186;48;5;186m▒\033[38;5;186;48;5;186m▒\033[38;5;220;48;5;185m▒\033[38;5;94;48;5;221m░\033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;186m▒\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;137m▒\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;101m▒\033[38;5;221;48;5;101m▒\033[38;5;94;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;137m▓\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;221m \033[38;5;172;48;5;221m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;180;48;5;95m▒\033[38;5;130;48;5;58m▒\033[38;5;179;48;5;58m░\033[38;5;94;48;5;58m▒\033[38;5;214;48;5;58m▒\033[38;5;179;48;5;58m▒\033[38;5;214;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;101m▒\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;180m▒\033[38;5;136;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;136;48;5;230m░\033[38;5;136;48;5;224m▒\033[38;5;220;48;5;223m▒\033[38;5;220;48;5;223m▒\033[38;5;220;48;5;223m░\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;186;48;5;186m▒\033[38;5;220;48;5;180m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;220;48;5;143m▒\033[38;5;178;48;5;179m▒\033[38;5;214;48;5;179m░\033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;136;48;5;180m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;101m▒\033[38;5;136;48;5;94m▒\033[38;5;221;48;5;58m░\033[38;5;179;48;5;95m▒\033[38;5;179;48;5;137m▓\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;214;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;221m \033[38;5;130;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;208;48;5;95m▒\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;58m░\033[38;5;179;48;5;58m▒\033[38;5;179;48;5;58m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;95m▒\033[38;5;94;48;5;95m▒\033[38;5;94;48;5;95m▓\033[38;5;214;48;5;144m▓\033[38;5;136;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;136;48;5;230m░\033[38;5;220;48;5;229m░\033[38;5;185;48;5;223m░\033[38;5;185;48;5;223m▒\033[38;5;185;48;5;187m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;220;48;5;186m▒\033[38;5;178;48;5;180m▒\033[38;5;178;48;5;180m▒\033[38;5;220;48;5;144m▒\033[38;5;178;48;5;144m▓\033[38;5;178;48;5;144m▓\033[38;5;178;48;5;186m▒\033[38;5;94;48;5;223m░\033[38;5;221;48;5;229m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;221;48;5;186m░\033[38;5;136;48;5;179m▒\033[38;5;178;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;221;48;5;137m▒\033[38;5;94;48;5;179m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;137;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;95m▒\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;94m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;95m▒\033[38;5;179;48;5;238m▒\033[38;5;179;48;5;240m▓\033[38;5;172;48;5;144m▓\033[38;5;220;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;144;48;5;253m▓\033[38;5;220;48;5;101m▓\033[38;5;187;48;5;150m▓\033[38;5;186;48;5;187m▒\033[38;5;143;48;5;144m▒\033[38;5;143;48;5;101m▓\033[38;5;144;48;5;143m▓\033[38;5;143;48;5;144m▓\033[38;5;187;48;5;180m▓\033[38;5;187;48;5;187m▒\033[38;5;185;48;5;193m▒\033[38;5;230;48;5;230m░\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;130;48;5;223m \033[38;5;130;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;222;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;137m▒\033[38;5;221;48;5;143m▒\033[38;5;221;48;5;179m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;180m▒\033[38;5;179;48;5;186m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;179;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;180;48;5;95m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;239m▒\033[38;5;172;48;5;239m▒\033[38;5;179;48;5;239m▒\033[38;5;179;48;5;240m▒\033[38;5;172;48;5;95m▓\033[38;5;172;48;5;137m▓\033[38;5;172;48;5;187m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;185;48;5;230m▒\033[38;5;187;48;5;254m▓\033[38;5;185;48;5;230m░\033[38;5;187;48;5;253m▓\033[38;5;144;48;5;187m▓\033[38;5;144;48;5;187m▓\033[38;5;186;48;5;255m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;220;48;5;229m \033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m░\033[38;5;172;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;94;48;5;143m▒\033[38;5;221;48;5;137m▒\033[38;5;136;48;5;137m▒\033[38;5;136;48;5;143m▒\033[38;5;136;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;172;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;131m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;238m▒\033[38;5;172;48;5;239m▒\033[38;5;172;48;5;239m▓\033[38;5;172;48;5;95m▓\033[38;5;172;48;5;101m▓\033[38;5;130;48;5;144m▓\033[38;5;223;48;5;224m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;220;48;5;229m \033[38;5;172;48;5;180m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;222;48;5;222m \033[38;5;214;48;5;221m \033[38;5;214;48;5;221m \033[38;5;172;48;5;221m░\033[38;5;179;48;5;179m░\033[38;5;214;48;5;179m▒\033[38;5;221;48;5;143m▒\033[38;5;178;48;5;137m▒\033[38;5;178;48;5;143m▒\033[38;5;178;48;5;143m▒\033[38;5;221;48;5;180m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;222m░\033[38;5;94;48;5;223m░\033[38;5;179;48;5;223m░\033[38;5;179;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;130;48;5;223m░\033[38;5;179;48;5;223m░\033[38;5;94;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;180;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;94m▒\033[38;5;179;48;5;58m░\033[38;5;94;48;5;58m▒\033[38;5;221;48;5;58m▒\033[38;5;179;48;5;237m▒\033[38;5;172;48;5;95m▓\033[38;5;172;48;5;181m▓\033[38;5;220;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;230m \033[38;5;178;48;5;223m░\033[38;5;221;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;214;48;5;221m \033[38;5;214;48;5;221m░\033[38;5;222;48;5;221m░\033[38;5;222;48;5;221m░\033[38;5;172;48;5;179m░\033[38;5;179;48;5;179m▒\033[38;5;214;48;5;143m▒\033[38;5;94;48;5;143m▒\033[38;5;94;48;5;180m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;223m░\033[38;5;94;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;222;48;5;223m░\033[38;5;179;48;5;223m░\033[38;5;214;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;179;48;5;222m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;208;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;58m▒\033[38;5;172;48;5;58m▒\033[38;5;130;48;5;101m▓\033[38;5;179;48;5;187m▒\033[38;5;220;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;136;48;5;229m░\033[38;5;221;48;5;223m░\033[38;5;136;48;5;186m▒\033[38;5;179;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;179m▒\033[38;5;179;48;5;179m▒\033[38;5;222;48;5;221m░\033[38;5;222;48;5;222m \033[38;5;214;48;5;222m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m░\033[38;5;94;48;5;186m░\033[38;5;214;48;5;186m░\033[38;5;172;48;5;223m░\033[38;5;130;48;5;181m▒\033[38;5;130;48;5;180m▒\033[38;5;172;48;5;181m▒\033[38;5;172;48;5;187m▒\033[38;5;172;48;5;223m░\033[38;5;222;48;5;224m \033[38;5;214;48;5;223m░\033[38;5;222;48;5;230m \033[38;5;222;48;5;230m \033[38;5;172;48;5;224m \033[38;5;172;48;5;224m \033[38;5;222;48;5;223m░\033[38;5;172;48;5;223m░\033[38;5;179;48;5;223m░\033[38;5;94;48;5;223m▒\033[38;5;221;48;5;187m▒\033[38;5;221;48;5;186m▒\033[38;5;178;48;5;180m▒\033[38;5;136;48;5;144m▒\033[38;5;221;48;5;143m▒\033[38;5;172;48;5;180m▒\033[38;5;130;48;5;216m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▓\033[38;5;137;48;5;137m▓\033[38;5;166;48;5;144m▓\033[38;5;166;48;5;188m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;136;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;178;48;5;187m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;186m▒\033[38;5;136;48;5;186m▒\033[38;5;94;48;5;186m▒\033[38;5;214;48;5;180m▒\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;186m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;223m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;178;48;5;230m \033[38;5;179;48;5;186m▒\033[38;5;130;48;5;180m▒\033[38;5;130;48;5;216m░\033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;137;48;5;137m▓\033[38;5;208;48;5;138m▓\033[38;5;178;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;231m \033[38;5;220;48;5;144m▓\033[38;5;220;48;5;101m▓\033[38;5;178;48;5;137m▓\033[38;5;221;48;5;179m▒\033[38;5;94;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;172;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m░\033[38;5;179;48;5;180m░\033[38;5;179;48;5;180m░\033[38;5;222;48;5;222m░\033[38;5;94;48;5;222m \033[38;5;136;48;5;222m \033[38;5;136;48;5;222m \033[38;5;178;48;5;222m \033[38;5;178;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;220;48;5;222m░\033[38;5;220;48;5;222m░\033[38;5;220;48;5;186m░\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;222;48;5;223m \033[38;5;130;48;5;222m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;209m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;180m▓\033[38;5;172;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;231m \033[38;5;94;48;5;187m▒\033[38;5;221;48;5;186m▒\033[38;5;221;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m░\033[38;5;214;48;5;222m░\033[38;5;222;48;5;222m \033[38;5;222;48;5;222m░\033[38;5;222;48;5;222m \033[38;5;214;48;5;222m \033[38;5;94;48;5;222m \033[38;5;221;48;5;222m \033[38;5;136;48;5;222m \033[38;5;178;48;5;222m \033[38;5;178;48;5;222m \033[38;5;178;48;5;222m \033[38;5;220;48;5;222m░\033[38;5;220;48;5;228m░\033[38;5;185;48;5;186m░\033[38;5;229;48;5;229m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;223m \033[38;5;130;48;5;222m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;137m▒\033[38;5;166;48;5;137m▒\033[38;5;214;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;230m \033[38;5;94;48;5;187m▒\033[38;5;221;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;222m░\033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;221;48;5;222m \033[38;5;221;48;5;222m \033[38;5;221;48;5;222m \033[38;5;136;48;5;222m \033[38;5;136;48;5;222m \033[38;5;178;48;5;222m░\033[38;5;220;48;5;222m░\033[38;5;229;48;5;229m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;178;48;5;229m \033[38;5;172;48;5;222m \033[38;5;172;48;5;221m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;220;48;5;230m \033[38;5;178;48;5;223m░\033[38;5;136;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;221;48;5;222m \033[38;5;221;48;5;222m \033[38;5;221;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;214;48;5;222m \033[38;5;222;48;5;222m \033[38;5;221;48;5;223m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;172;48;5;223m \033[38;5;130;48;5;222m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;221;48;5;224m░\033[38;5;220;48;5;187m▒\033[38;5;178;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;178;48;5;222m░\033[38;5;136;48;5;186m▒\033[38;5;136;48;5;179m▒\033[38;5;136;48;5;186m▒\033[38;5;178;48;5;222m░\033[38;5;136;48;5;222m░\033[38;5;94;48;5;223m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;172;48;5;223m \033[38;5;130;48;5;216m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;172;48;5;222m \033[38;5;130;48;5;216m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;166;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;220;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;229m \033[38;5;130;48;5;222m \033[38;5;130;48;5;216m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;215;48;5;215m \033[38;5;166;48;5;215m░\033[38;5;166;48;5;215m░\033[38;5;166;48;5;173m░\033[38;5;166;48;5;173m▒\033[38;5;180;48;5;181m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;94;48;5;223m \033[38;5;172;48;5;222m \033[38;5;130;48;5;216m \033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;208;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;215;48;5;215m░\033[38;5;180;48;5;173m▒\033[38;5;166;48;5;180m▒\033[38;5;94;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;94;48;5;223m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;215;48;5;215m░\033[38;5;180;48;5;179m▒\033[38;5;166;48;5;216m░\033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;230;48;5;230m \033[38;5;214;48;5;223m░\033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;222m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m \033[38;5;215;48;5;215m \033[38;5;208;48;5;179m░\033[38;5;180;48;5;179m▒\033[38;5;166;48;5;223m░\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m░\033[38;5;94;48;5;187m▒\033[38;5;172;48;5;186m▒\033[38;5;172;48;5;222m░\033[38;5;130;48;5;222m░\033[38;5;130;48;5;222m \033[38;5;172;48;5;222m \033[38;5;130;48;5;215m \033[38;5;166;48;5;215m \033[38;5;215;48;5;179m░\033[38;5;180;48;5;173m▒\033[38;5;180;48;5;173m▒\033[38;5;172;48;5;224m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;181m▓\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;180m▒\033[38;5;172;48;5;216m░\033[38;5;172;48;5;180m░\033[38;5;130;48;5;179m░\033[38;5;130;48;5;179m░\033[38;5;130;48;5;179m▒\033[38;5;130;48;5;179m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;180m▒\033[38;5;94;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");
    		$display("\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;144m▓\033[38;5;172;48;5;101m▓\033[38;5;172;48;5;144m▓\033[38;5;214;48;5;137m▓\033[38;5;94;48;5;143m▒\033[38;5;179;48;5;180m▒\033[38;5;94;48;5;143m▓\033[38;5;178;48;5;95m▓\033[38;5;220;48;5;137m▓\033[38;5;220;48;5;223m▒\033[38;5;230;48;5;230m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[0m");

			$display("\nThere is some bug in your code. Errors exceed 100.\n");
			$finish;
		end
	end

endmodule





