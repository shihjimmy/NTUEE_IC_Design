`timescale 1ns / 1ps
`define CYCLE 7.8
`define PATTERN 1000

module tb;

//clk generation
reg clk = 1;
always #(`CYCLE/2) clk = ~clk;

//dump waveform
initial begin
	$fsdbDumpfile("factor.fsdb");
	$fsdbDumpvars(0,"+mda");
end

//time out
initial begin
	#(100000*`CYCLE);
	FAIL;
	$display("\n\033[1;31m=============================================");
	$display("           Simulation Time Out!      ");
	$display("=============================================\033[0m");
	$finish;
end

//instatiate DUT
reg rst_n = 1;
reg [11:0] n;
reg in_valid;
wire out_valid;
wire [3:0] p2;
wire [2:0] p3;
wire [2:0] p5;
wire [50:0] number;

factor DUT(
	.clk(clk),
	.rst_n(rst_n),
	.i_n(n),
	.i_in_valid(in_valid),
	.o_out_valid(out_valid),
	.o_p2(p2),
	.o_p3(p3),
	.o_p5(p5),
	.number(number)
);

//Initial memory
reg [12:0] INPUT_N_MEM [0:`PATTERN-1];
reg [3:0]  GOLDEN_2_MEM [0:`PATTERN-1];
reg [2:0]  GOLDEN_3_MEM [0:`PATTERN-1];
reg [2:0]  GOLDEN_5_MEM [0:`PATTERN-1];

initial begin
	$readmemb("pattern/Inn.dat",  INPUT_N_MEM);
	$readmemb("pattern/Gol2.dat", GOLDEN_2_MEM);
	$readmemb("pattern/Gol3.dat", GOLDEN_3_MEM);
	$readmemb("pattern/Gol5.dat", GOLDEN_5_MEM);
end

//Latency
integer latency;
`ifdef PIPELINE
	always @(posedge clk or negedge rst_n) begin 
		if (~rst_n) begin 
			latency = -1;
		end
		else begin
			latency = latency + 1;
		end
	end
`else
	always @(posedge clk or negedge rst_n) begin 
		if (~rst_n) begin 
			latency = -1;
		end
		else begin
			latency = latency + 1;
		end
	end
`endif

//input pattern & check result
integer i,j;
integer err_num = 0;
integer total_latency = 0;

`ifdef PIPELINE
//input
initial begin
	//reset 
	in_valid = 0;
	@(posedge clk) rst_n = 0;
	@(posedge clk); 
	rst_n = 1;
	@(posedge clk);
	for (i=0; i<`PATTERN; i=i+1) begin
		#(0.6); //filp flop hold time
		n = INPUT_N_MEM[i];
		in_valid = 1;
		@(posedge clk); 
	end
	#(0.6);
	in_valid = 0;
	n = 'bx;
end

//check output
initial begin
	wait (out_valid);
	@(negedge clk);
	for (j=0; j<`PATTERN; j=j+1) begin
		if (out_valid !== 1)begin
			FAIL;
			$display("\n\033[1;31m=============================================");
			$display("     out_valid should be kept high once      ");
			$display("     you pull it up in pipeline mode.       ");
			$display("=============================================\033[0m");
			@(negedge clk);
			$finish;
		end else if (GOLDEN_2_MEM[j] === p2 && GOLDEN_3_MEM[j] === p3 && GOLDEN_5_MEM[j] === p5 && p2!==4'bx && p3 !== 3'bx && p5 !== 3'bx) begin
			`ifdef DEBUG
				$display("\033[1;92mPattern %3d passed. / Input N:%4d / Output P2:%2d / Output P3: %1d / Output P5: %1d / Golden P2: %1d / Golden P3: %1d/ Golden P5: %1d\033[0m", j, INPUT_N_MEM[j], p2, p3, p5, GOLDEN_2_MEM[j], GOLDEN_3_MEM[j], GOLDEN_5_MEM[j]);
			`endif
		end else begin
			`ifdef DEBUG
				$display("\033[1;31mPattern %3d failed. / Input N:%4d / Output P2:%2d / Output P3: %1d / Output P5: %1d / Golden P2: %1d / Golden P3: %1d/ Golden P5: %1d\033[0m", j, INPUT_N_MEM[j], p2, p3, p5, GOLDEN_2_MEM[j], GOLDEN_3_MEM[j], GOLDEN_5_MEM[j]);
			`endif
			err_num = err_num + 1;
		end
		@(negedge clk);
	end
	total_latency = latency-1;

	if (err_num != 0) begin
		FAIL;
		$display("\n\033[1;31m=============================================");
		$display("              Simulation failed              ");
		$display("=============================================\033[0m");
	end
	else begin
		PASS;
		$display("\n\033[1;92m=============================================");
		$display("              Simulation passed              ");
		$display("=============================================\033[0m");
	end

	$display("\n\033[1;96m=============================================");
	$display("                   Summary                   ");
	$display("=============================================");
	$display("  	Clock cycle:           %.1f ns", `CYCLE);
	$display("  	Number of transistors: %.0f", $itor(number));
	$display("  	Total excution cycle:  %.0f", $itor(total_latency));
	$display("  	Correctness Score:     %.1f", 40.0 * $itor($itor(`PATTERN) - $itor(err_num)) / $itor(`PATTERN));
	$display("  	Performance Score:     %.1f", $itor(total_latency) * $itor(number) * `CYCLE);
	$display("=============================================\033[0m");

	$finish;
end

`else 
initial begin
	in_valid = 0;
	rst_n = 1;
	@(posedge clk)
	for (i=0; i<`PATTERN; i=i+1) begin
		//reset 
		rst_n = 0;
		@(posedge clk); 
		rst_n = 1;
		@(posedge clk);
		#(0.6); //filp flop hold time
		in_valid = 1;
		n = INPUT_N_MEM[i];

		wait (out_valid);
		@(negedge clk);
		j=i;
		total_latency = total_latency + latency;
		if (GOLDEN_2_MEM[j] === p2 && GOLDEN_3_MEM[j] === p3 && GOLDEN_5_MEM[j] === p5 && p2!==4'bx && p3 !== 3'bx && p5 !== 3'bx) begin
			`ifdef DEBUG
				$display("\033[1;92mPattern %3d passed. / Input N:%4d / Output P2:%2d / Output P3: %1d / Output P5: %1d / Golden P2: %1d / Golden P3: %1d/ Golden P5: %1d\033[0m", j, INPUT_N_MEM[j], p2, p3, p5, GOLDEN_2_MEM[j], GOLDEN_3_MEM[j], GOLDEN_5_MEM[j]);
			`endif
		end
		else begin
			`ifdef DEBUG
				$display("\033[1;31mPattern %3d failed. / Input N:%4d / Output P2:%2d / Output P3: %1d / Output P5: %1d / Golden P2: %1d / Golden P3: %1d/ Golden P5: %1d\033[0m", j, INPUT_N_MEM[j], p2, p3, p5, GOLDEN_2_MEM[j], GOLDEN_3_MEM[j], GOLDEN_5_MEM[j]);
			`endif
			err_num = err_num + 1;
		end
		@(posedge clk);
		n = 'bx;
		in_valid = 0;
	end

	if (err_num != 0) begin
		FAIL;
		$display("\n\033[1;31m=============================================");
		$display("              Simulation failed              ");
		$display("=============================================\033[0m");
	end
	else begin 
		PASS;
		$display("\n\033[1;92m=============================================");
		$display("              Simulation passed              ");
		$display("=============================================\033[0m");
	end

	$display("\n\033[1;96m=============================================");
	$display("                   Summary                   ");
	$display("=============================================");
	$display("  	Clock cycle:           %.1f ns", `CYCLE);
	$display("  	Number of transistors: %.0f", $itor(number));
	$display("  	Total excution cycle:  %.0f", $itor(total_latency));
	$display("  	Correctness Score:     %.1f", 40.0 * $itor($itor(`PATTERN) - $itor(err_num)) / $itor(`PATTERN));
	$display("  	Performance Score:     %.1f", $itor(total_latency) * $itor(number) * `CYCLE);
	$display("=============================================\033[0m");

	@(negedge clk);
	$finish;
end
`endif

task PASS;
begin
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[38;5;204;48;5;232m \033[38;5;126;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;89;48;5;22m░\033[38;5;212;48;5;22m░\033[38;5;204;48;5;16m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;204;48;5;232m \033[38;5;126;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;126;48;5;22m░\033[38;5;204;48;5;232m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;161;48;5;233m░\033[38;5;212;48;5;22m░\033[38;5;126;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;89;48;5;22m░\033[38;5;162;48;5;22m░\033[38;5;204;48;5;16m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;125;48;5;22m░\033[38;5;199;48;5;22m░\033[38;5;126;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;163;48;5;22m░\033[38;5;126;48;5;22m░\033[38;5;199;48;5;22m░\033[38;5;125;48;5;22m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;52;48;5;232m░\033[38;5;98;48;5;235m▒\033[38;5;61;48;5;235m▓\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;84;48;5;173m░\033[38;5;41;48;5;209m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[38;5;212;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;62;48;5;41m░\033[38;5;92;48;5;2m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;99;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;176;48;5;41m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;125;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;212;48;5;41m░\033[0m \033[0m \033[0m \033[38;5;56;48;5;41m░\033[38;5;99;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;56;48;5;2m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;208;48;5;236m▓\033[38;5;95;48;5;234m▓\033[38;5;166;48;5;237m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;84;48;5;208m▒\033[38;5;222;48;5;223m \033[38;5;166;48;5;209m \033[38;5;190;48;5;208m▓\033[38;5;41;48;5;209m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;238m▓\033[38;5;85;48;5;208m░\033[38;5;85;48;5;208m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[38;5;212;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;57;48;5;2m░\033[38;5;125;48;5;22m░\033[38;5;165;48;5;22m░\033[38;5;99;48;5;41m░\033[38;5;56;48;5;41m▒\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;141;48;5;34m░\033[0m \033[0m \033[0m \033[38;5;57;48;5;35m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;99;48;5;41m▒\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;99;48;5;35m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;53;48;5;22m░\033[38;5;62;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;62;48;5;41m░\033[38;5;99;48;5;41m░\033[38;5;92;48;5;28m░\033[38;5;125;48;5;22m░\033[38;5;57;48;5;41m░\033[38;5;99;48;5;41m░\033[38;5;20;48;5;41m░\033[38;5;20;48;5;41m░\033[0m \033[0m \033[38;5;141;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;126;48;5;41m▒\033[38;5;99;48;5;41m░\033[38;5;125;48;5;22m░\033[38;5;162;48;5;22m░\033[38;5;99;48;5;41m░\033[38;5;99;48;5;41m░\033[38;5;134;48;5;41m▒\033[38;5;135;48;5;2m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;190;48;5;235m░\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;179m░\033[38;5;95;48;5;235m▓\033[38;5;220;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;49;48;5;222m░\033[38;5;67;48;5;208m▒\033[38;5;136;48;5;222m \033[38;5;172;48;5;221m \033[38;5;41;48;5;209m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;166;48;5;235m▒\033[38;5;85;48;5;208m░\033[38;5;223;48;5;222m \033[38;5;230;48;5;231m \033[38;5;166;48;5;216m \033[38;5;84;48;5;209m▒\033[38;5;85;48;5;208m░\033[38;5;76;48;5;95m▓\033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[38;5;212;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;165;48;5;22m░\033[0m \033[0m \033[0m \033[38;5;55;48;5;41m \033[38;5;84;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;19;48;5;34m░\033[0m \033[0m \033[38;5;177;48;5;34m░\033[38;5;99;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;20;48;5;41m░\033[38;5;135;48;5;41m░\033[38;5;84;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;55;48;5;28m░\033[0m \033[0m \033[0m \033[0m \033[38;5;53;48;5;22m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;20;48;5;41m░\033[38;5;204;48;5;232m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;99;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;135;48;5;28m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;167;48;5;233m░\033[38;5;42;48;5;235m▒\033[38;5;95;48;5;235m▓\033[38;5;130;48;5;95m▒\033[38;5;222;48;5;222m \033[38;5;221;48;5;222m \033[38;5;172;48;5;179m░\033[38;5;209;48;5;235m▓\033[38;5;65;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;115;48;5;137m▒\033[38;5;41;48;5;209m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;173;48;5;240m▓\033[38;5;71;48;5;94m▓\033[38;5;85;48;5;209m░\033[38;5;35;48;5;208m▒\033[38;5;136;48;5;222m \033[38;5;130;48;5;215m \033[38;5;85;48;5;209m░\033[38;5;209;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[38;5;212;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;165;48;5;22m░\033[0m \033[38;5;204;48;5;16m \033[38;5;204;48;5;232m░\033[38;5;99;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;57;48;5;28m░\033[0m \033[38;5;204;48;5;16m \033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;99;48;5;34m░\033[38;5;204;48;5;16m \033[38;5;141;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;99;48;5;41m▒\033[0m \033[0m \033[0m \033[0m \033[38;5;200;48;5;22m \033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;20;48;5;41m░\033[38;5;57;48;5;35m░\033[38;5;204;48;5;16m \033[0m \033[0m \033[0m \033[0m \033[38;5;56;48;5;41m░\033[38;5;21;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;62;48;5;41m░\033[38;5;99;48;5;41m░\033[38;5;204;48;5;232m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;137;48;5;235m▓\033[38;5;75;48;5;234m░\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;172;48;5;137m▒\033[38;5;214;48;5;221m \033[38;5;172;48;5;215m \033[38;5;130;48;5;173m▒\033[38;5;209;48;5;235m▓\033[38;5;65;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;209;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;233m░\033[38;5;85;48;5;208m░\033[38;5;85;48;5;208m░\033[38;5;209;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[38;5;212;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;99;48;5;41m░\033[38;5;55;48;5;28m░\033[0m \033[38;5;204;48;5;16m \033[38;5;141;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;134;48;5;41m▒\033[0m \033[0m \033[38;5;197;48;5;233m \033[38;5;165;48;5;41m▒\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;19;48;5;35m░\033[0m \033[0m \033[0m \033[0m \033[38;5;204;48;5;16m \033[38;5;55;48;5;35m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;62;48;5;41m░\033[38;5;56;48;5;34m░\033[0m \033[0m \033[0m \033[38;5;198;48;5;22m \033[38;5;141;48;5;41m░\033[38;5;176;48;5;41m▒\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;205;48;5;41m░\033[38;5;206;48;5;22m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;173;48;5;234m▓\033[38;5;119;48;5;235m░\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;95m▓\033[38;5;94;48;5;186m░\033[38;5;222;48;5;222m░\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;94m▒\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;234m▒\033[38;5;197;48;5;235m░\033[38;5;209;48;5;235m▓\033[38;5;197;48;5;235m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[38;5;212;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;98;48;5;41m▒\033[38;5;200;48;5;41m▒\033[38;5;163;48;5;41m▒\033[38;5;20;48;5;41m░\033[38;5;99;48;5;41m░\033[38;5;55;48;5;28m░\033[38;5;204;48;5;232m \033[0m \033[0m \033[0m \033[38;5;56;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;21;48;5;41m░\033[38;5;140;48;5;41m▒\033[38;5;140;48;5;41m▒\033[38;5;140;48;5;41m▒\033[38;5;99;48;5;41m▒\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;57;48;5;41m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;125;48;5;22m \033[38;5;171;48;5;2m░\033[38;5;99;48;5;41m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;177;48;5;22m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;5;48;5;2m░\033[38;5;135;48;5;34m░\033[38;5;125;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;99;48;5;41m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;166;48;5;236m▓\033[38;5;42;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;237m▓\033[38;5;172;48;5;101m▒\033[38;5;179;48;5;179m░\033[38;5;136;48;5;222m \033[38;5;179;48;5;179m░\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;166;48;5;236m▒\033[38;5;119;48;5;235m░\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;52;48;5;232m░\033[38;5;119;48;5;236m▓\033[38;5;82;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;238m▓\033[38;5;208;48;5;58m▒\033[38;5;209;48;5;235m▓\033[38;5;113;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;107;48;5;94m▓\033[38;5;114;48;5;208m▒\033[38;5;41;48;5;172m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[38;5;212;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;165;48;5;22m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;161;48;5;233m░\033[38;5;56;48;5;41m▒\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;20;48;5;41m░\033[38;5;204;48;5;232m \033[0m \033[38;5;200;48;5;22m░\033[38;5;99;48;5;41m░\033[38;5;204;48;5;16m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;135;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;93;48;5;22m░\033[0m \033[38;5;57;48;5;41m░\033[38;5;135;48;5;41m░\033[38;5;204;48;5;16m \033[0m \033[0m \033[0m \033[0m \033[38;5;204;48;5;232m \033[38;5;99;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;202;48;5;236m▓\033[38;5;204;48;5;235m▒\033[38;5;95;48;5;234m▓\033[38;5;166;48;5;236m▓\033[38;5;172;48;5;95m▓\033[38;5;222;48;5;222m░\033[38;5;136;48;5;222m \033[38;5;94;48;5;221m \033[38;5;222;48;5;215m \033[38;5;172;48;5;137m▒\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;179m░\033[38;5;94;48;5;221m \033[38;5;172;48;5;137m▒\033[38;5;172;48;5;131m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;94m▒\033[38;5;204;48;5;234m▓\033[38;5;179;48;5;236m▓\033[0m \033[38;5;173;48;5;236m▓\033[38;5;84;48;5;236m▓\033[38;5;119;48;5;235m░\033[38;5;204;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;240m▓\033[38;5;179;48;5;179m▒\033[38;5;94;48;5;222m \033[38;5;221;48;5;222m \033[38;5;130;48;5;173m░\033[38;5;204;48;5;234m▓\033[38;5;72;48;5;235m▓\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;41;48;5;209m░\033[38;5;208;48;5;216m \033[38;5;94;48;5;230m \033[38;5;166;48;5;208m░\033[38;5;41;48;5;208m░\033[38;5;209;48;5;234m░\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[38;5;212;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;165;48;5;22m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;161;48;5;22m \033[38;5;99;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;20;48;5;41m░\033[38;5;53;48;5;22m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;165;48;5;2m░\033[38;5;99;48;5;41m▒\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;125;48;5;41m░\033[0m \033[38;5;53;48;5;22m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;20;48;5;41m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;99;48;5;41m░\033[38;5;200;48;5;22m░\033[0m \033[38;5;99;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;20;48;5;41m░\033[38;5;20;48;5;41m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;99;48;5;41m░\033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;119;48;5;235m▓\033[38;5;119;48;5;235m░\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;239m▓\033[38;5;179;48;5;137m▒\033[38;5;222;48;5;222m░\033[38;5;214;48;5;222m \033[38;5;214;48;5;221m \033[38;5;214;48;5;221m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;173m▒\033[38;5;222;48;5;215m \033[38;5;94;48;5;221m \033[38;5;172;48;5;179m░\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;137m▒\033[38;5;138;48;5;234m▓\033[38;5;208;48;5;238m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;137m▒\033[38;5;179;48;5;179m▒\033[38;5;222;48;5;222m░\033[38;5;179;48;5;215m░\033[38;5;172;48;5;137m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;179m▒\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;136m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;202;48;5;236m▓\033[38;5;137;48;5;237m▒\033[38;5;202;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;61;48;5;235m▓\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;113;48;5;94m▓\033[38;5;178;48;5;208m▒\033[38;5;208;48;5;222m \033[38;5;230;48;5;230m \033[38;5;229;48;5;229m \033[38;5;229;48;5;229m \033[38;5;230;48;5;230m \033[38;5;166;48;5;209m \033[38;5;48;48;5;208m░\033[38;5;190;48;5;95m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[38;5;212;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;165;48;5;22m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;141;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;57;48;5;34m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;141;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;135;48;5;2m░\033[38;5;200;48;5;22m░\033[38;5;20;48;5;41m░\033[38;5;62;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;62;48;5;41m░\033[38;5;20;48;5;41m░\033[38;5;92;48;5;28m░\033[0m \033[0m \033[0m \033[38;5;57;48;5;41m░\033[38;5;171;48;5;41m▒\033[38;5;20;48;5;41m░\033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;84;48;5;41m \033[38;5;99;48;5;41m▒\033[38;5;99;48;5;35m░\033[38;5;171;48;5;237m▒\033[38;5;41;48;5;236m▓\033[38;5;55;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;222m░\033[38;5;94;48;5;221m \033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;179m░\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;173m▒\033[38;5;173;48;5;235m▓\033[38;5;180;48;5;238m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;95m▒\033[38;5;172;48;5;173m░\033[38;5;130;48;5;173m░\033[38;5;208;48;5;238m▒\033[38;5;173;48;5;235m▓\033[38;5;172;48;5;137m▒\033[38;5;94;48;5;221m \033[38;5;222;48;5;215m \033[38;5;94;48;5;221m \033[38;5;172;48;5;95m▒\033[38;5;95;48;5;235m▓\033[38;5;204;48;5;95m▓\033[38;5;204;48;5;138m▒\033[38;5;204;48;5;95m▓\033[38;5;209;48;5;234m▓\033[38;5;78;48;5;236m▓\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;220;48;5;58m▓\033[38;5;48;48;5;209m░\033[38;5;166;48;5;209m░\033[38;5;178;48;5;222m \033[38;5;228;48;5;228m \033[38;5;166;48;5;208m░\033[38;5;71;48;5;130m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;172;48;5;236m▓\033[38;5;55;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;234m▓\033[38;5;130;48;5;95m▒\033[38;5;221;48;5;222m \033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;173m▒\033[38;5;202;48;5;235m▓\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;179m░\033[38;5;172;48;5;179m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;137m▒\033[38;5;166;48;5;237m▒\033[38;5;204;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;236m▓\033[38;5;197;48;5;234m▓\033[38;5;197;48;5;234m▓\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;174m▒\033[38;5;204;48;5;174m▒\033[38;5;197;48;5;211m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;52;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;41;48;5;208m░\033[38;5;166;48;5;208m░\033[38;5;41;48;5;209m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;244m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;197;48;5;235m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;173m▒\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;137m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;221m░\033[38;5;94;48;5;222m \033[38;5;214;48;5;221m \033[38;5;179;48;5;179m░\033[38;5;172;48;5;215m░\033[38;5;222;48;5;221m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;95m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;236m▓\033[38;5;168;48;5;175m▒\033[38;5;204;48;5;175m░\033[38;5;211;48;5;211m░\033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;204;48;5;131m▓\033[38;5;173;48;5;235m▓\033[38;5;41;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;66;48;5;244m▓\033[38;5;209;48;5;234m▓\033[38;5;133;48;5;235m▓\033[38;5;40;48;5;235m░\033[38;5;95;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;95;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;236m▓\033[38;5;172;48;5;137m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;130;48;5;173m░\033[38;5;130;48;5;94m▒\033[38;5;173;48;5;235m▓\033[38;5;166;48;5;237m▒\033[38;5;130;48;5;136m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;137m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;204;48;5;237m▓\033[38;5;197;48;5;175m▒\033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;52;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;41;48;5;209m░\033[38;5;119;48;5;208m▒\033[38;5;76;48;5;94m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;138;48;5;238m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;236m▓\033[38;5;166;48;5;237m▒\033[38;5;172;48;5;215m░\033[38;5;94;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;166;48;5;236m▒\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;234m▓\033[38;5;130;48;5;131m▒\033[38;5;94;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;180;48;5;237m▒\033[38;5;137;48;5;237m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;215m \033[38;5;214;48;5;221m \033[38;5;172;48;5;179m░\033[38;5;137;48;5;237m▒\033[38;5;180;48;5;238m▒\033[38;5;172;48;5;131m▒\033[38;5;130;48;5;179m░\033[38;5;130;48;5;215m \033[38;5;130;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;166;48;5;237m▒\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;168;48;5;175m▒\033[38;5;218;48;5;218m \033[38;5;204;48;5;95m▓\033[38;5;209;48;5;235m▓\033[38;5;191;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;173;48;5;234m▒\033[38;5;166;48;5;208m░\033[38;5;230;48;5;230m \033[38;5;208;48;5;222m \033[38;5;41;48;5;208m░\033[38;5;85;48;5;208m░\033[38;5;71;48;5;130m▓\033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;173;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;95m▓\033[38;5;204;48;5;211m░\033[38;5;204;48;5;174m▒\033[38;5;95;48;5;238m▓\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;166;48;5;236m▓\033[38;5;95;48;5;235m▓\033[38;5;166;48;5;236m▓\033[38;5;172;48;5;179m░\033[38;5;214;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;221m \033[38;5;172;48;5;179m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;179m░\033[38;5;130;48;5;173m▒\033[38;5;172;48;5;173m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;166;48;5;237m▒\033[38;5;209;48;5;234m▓\033[38;5;138;48;5;236m▓\033[38;5;168;48;5;138m▒\033[38;5;173;48;5;235m▓\033[38;5;197;48;5;235m░\033[0m \033[0m \033[0m \033[0m \033[38;5;42;48;5;138m▓\033[38;5;80;48;5;209m▒\033[38;5;166;48;5;215m░\033[38;5;209;48;5;208m \033[38;5;84;48;5;130m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;191;48;5;240m▓\033[38;5;41;48;5;208m░\033[38;5;215;48;5;208m░\033[38;5;228;48;5;228m \033[38;5;228;48;5;228m \033[38;5;166;48;5;209m░\033[38;5;84;48;5;130m▒\033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;234m▒\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;95m▓\033[38;5;204;48;5;211m░\033[38;5;204;48;5;174m▒\033[38;5;204;48;5;174m▒\033[38;5;204;48;5;211m░\033[38;5;204;48;5;95m▓\033[38;5;166;48;5;236m▒\033[38;5;172;48;5;179m░\033[38;5;208;48;5;58m▒\033[38;5;95;48;5;235m▓\033[38;5;202;48;5;235m▓\033[38;5;172;48;5;173m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;179m░\033[38;5;137;48;5;237m▒\033[38;5;180;48;5;58m▒\033[38;5;130;48;5;173m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;179m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;133;48;5;235m▓\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[38;5;85;48;5;209m░\033[38;5;84;48;5;208m░\033[38;5;222;48;5;221m \033[38;5;84;48;5;208m▒\033[38;5;136;48;5;58m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;41;48;5;208m░\033[38;5;166;48;5;208m░\033[38;5;85;48;5;209m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;149;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;95m▓\033[38;5;218;48;5;218m \033[38;5;204;48;5;211m░\033[38;5;204;48;5;174m▒\033[38;5;204;48;5;174m▒\033[38;5;204;48;5;175m░\033[38;5;204;48;5;174m▒\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;234m▓\033[38;5;172;48;5;137m▒\033[38;5;214;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;179m░\033[38;5;166;48;5;236m▓\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;231;48;5;231m▓\033[38;5;178;48;5;230m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;173m░\033[38;5;130;48;5;94m▒\033[38;5;166;48;5;237m▒\033[38;5;172;48;5;179m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;221m \033[38;5;208;48;5;238m▒\033[38;5;209;48;5;235m▓\033[38;5;99;48;5;235m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;78;48;5;173m▒\033[38;5;154;48;5;94m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;149;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;95m▓\033[38;5;218;48;5;218m \033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;211;48;5;211m░\033[38;5;204;48;5;95m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;94;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;229m \033[38;5;222;48;5;221m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;221m \033[38;5;172;48;5;95m▒\033[38;5;137;48;5;237m▒\033[38;5;208;48;5;237m▒\033[38;5;208;48;5;237m▒\033[38;5;137;48;5;237m▒\033[38;5;137;48;5;237m▒\033[38;5;166;48;5;236m▓\033[38;5;202;48;5;236m▓\033[38;5;173;48;5;235m▓\033[38;5;166;48;5;237m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;221m \033[38;5;172;48;5;137m▒\033[38;5;95;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;234m▒\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;240m▓\033[38;5;218;48;5;218m \033[38;5;161;48;5;218m \033[38;5;218;48;5;218m \033[38;5;204;48;5;95m▓\033[38;5;209;48;5;234m▓\033[38;5;166;48;5;236m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;229m \033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;130m░\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;238m▓\033[38;5;218;48;5;218m \033[38;5;218;48;5;218m \033[38;5;204;48;5;95m▓\033[38;5;209;48;5;234m▓\033[38;5;166;48;5;236m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;137m▒\033[38;5;180;48;5;237m▒\033[38;5;202;48;5;236m▓\033[38;5;172;48;5;179m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;231m▒\033[38;5;181;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;230m \033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;130m░\033[38;5;95;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;236m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;209;48;5;235m▓\033[38;5;138;48;5;237m▓\033[38;5;218;48;5;218m \033[38;5;204;48;5;132m▓\033[38;5;173;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;221m \033[38;5;214;48;5;221m \033[38;5;94;48;5;221m \033[38;5;222;48;5;215m \033[38;5;172;48;5;179m░\033[38;5;172;48;5;137m▒\033[38;5;180;48;5;238m▒\033[38;5;173;48;5;235m▓\033[38;5;137;48;5;237m▒\033[38;5;130;48;5;130m▒\033[38;5;172;48;5;179m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;209;48;5;252m▓\033[38;5;209;48;5;242m▓\033[38;5;173;48;5;237m▓\033[38;5;209;48;5;237m▓\033[38;5;209;48;5;59m▓\033[38;5;209;48;5;240m▓\033[38;5;209;48;5;234m▓\033[38;5;173;48;5;234m▓\033[38;5;209;48;5;234m▓\033[38;5;173;48;5;237m▓\033[38;5;209;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;138;48;5;231m▓\033[38;5;173;48;5;248m▓\033[38;5;173;48;5;235m▓\033[38;5;173;48;5;244m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;94;48;5;222m \033[38;5;222;48;5;221m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;208;48;5;94m░\033[38;5;95;48;5;235m▓\033[38;5;133;48;5;235m▓\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;55;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;168;48;5;175m▒\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;234m▓\033[38;5;172;48;5;173m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;173m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;209;48;5;245m▓\033[38;5;209;48;5;236m▓\033[38;5;137;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;202;48;5;253m▓\033[38;5;173;48;5;102m▓\033[38;5;173;48;5;236m▓\033[38;5;209;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;245m▓\033[38;5;209;48;5;242m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;229m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;202;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;191;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;202;48;5;234m▓\033[38;5;42;48;5;235m▒\033[38;5;197;48;5;235m░\033[38;5;35;48;5;236m▓\033[38;5;167;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;175;48;5;235m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;178;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;249;48;5;249m▓\033[38;5;209;48;5;238m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;247m▓\033[38;5;209;48;5;242m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;253m▓\033[38;5;173;48;5;238m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;229m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;137m▒\033[38;5;204;48;5;234m▓\033[38;5;129;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;79;48;5;236m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;173;48;5;247m▓\033[38;5;218;48;5;218m \033[38;5;161;48;5;224m \033[38;5;249;48;5;249m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;137;48;5;236m▓\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;190;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;202;48;5;253m▓\033[38;5;209;48;5;236m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;173;48;5;235m▓\033[38;5;173;48;5;234m▓\033[38;5;166;48;5;244m▓\033[38;5;222;48;5;231m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;136;48;5;231m \033[38;5;166;48;5;248m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;214m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;80;48;5;251m▒\033[38;5;1;48;5;233m░\033[38;5;79;48;5;236m▒\033[38;5;173;48;5;234m▓\033[38;5;209;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;239m▓\033[38;5;209;48;5;59m▓\033[38;5;168;48;5;7m▓\033[38;5;197;48;5;175m░\033[38;5;197;48;5;218m░\033[38;5;209;48;5;249m▓\033[38;5;209;48;5;237m▓\033[38;5;53;48;5;235m░\033[38;5;209;48;5;234m▒\033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;199;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;253m▓\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;243m▓\033[38;5;166;48;5;188m▒\033[38;5;166;48;5;255m░\033[38;5;223;48;5;230m░\033[38;5;202;48;5;188m▓\033[38;5;166;48;5;102m▓\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;138m▒\033[38;5;204;48;5;211m░\033[38;5;204;48;5;174m▒\033[38;5;204;48;5;239m▓\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;238m▓\033[38;5;209;48;5;239m▓\033[38;5;209;48;5;102m▓\033[38;5;180;48;5;255m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;166;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;84;48;5;236m▓\033[38;5;46;48;5;235m░\033[38;5;173;48;5;236m▓\033[38;5;209;48;5;255m▓\033[38;5;225;48;5;231m \033[38;5;197;48;5;211m░\033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;125;48;5;225m \033[38;5;231;48;5;231m▓\033[38;5;216;48;5;231m \033[38;5;209;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;61;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;52;48;5;232m░\033[38;5;104;48;5;235m▒\033[38;5;204;48;5;234m▓\033[38;5;172;48;5;173m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;254m▓\033[38;5;137;48;5;250m▓\033[38;5;166;48;5;145m▓\033[38;5;137;48;5;187m▓\033[38;5;230;48;5;231m \033[38;5;209;48;5;237m▓\033[38;5;197;48;5;211m░\033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;204;48;5;132m▓\033[38;5;173;48;5;241m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;172m░\033[38;5;166;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;126;48;5;225m \033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;163;48;5;225m \033[38;5;231;48;5;231m▓\033[38;5;125;48;5;224m \033[38;5;161;48;5;218m \033[38;5;225;48;5;231m \033[38;5;209;48;5;250m▓\033[38;5;209;48;5;234m▓\033[38;5;110;48;5;235m▒\033[0m░\033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;251m▓\033[38;5;95;48;5;238m▓\033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;204;48;5;95m▓\033[38;5;173;48;5;102m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;237m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;223;48;5;230m \033[38;5;173;48;5;247m▓\033[38;5;209;48;5;234m▓\033[38;5;133;48;5;235m▓\033[38;5;1;48;5;232m░\033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;94;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;247m▓\033[38;5;204;48;5;238m▓\033[38;5;204;48;5;95m▓\033[38;5;209;48;5;237m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;130m░\033[38;5;204;48;5;234m▓\033[38;5;95;48;5;234m▓\033[38;5;172;48;5;179m░\033[38;5;214;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;223;48;5;231m \033[38;5;166;48;5;224m░\033[38;5;137;48;5;145m▓\033[38;5;173;48;5;237m▓\033[38;5;173;48;5;235m▓\033[38;5;211;48;5;235m░\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;243;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;119;48;5;238m▓\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;236m▓\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;221m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;166;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;214;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;102m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;133;48;5;235m▓\033[38;5;220;48;5;235m▓\033[38;5;88;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;235m▓\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;223m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;94m▒\033[38;5;204;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;172;48;5;221m \033[38;5;130;48;5;95m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;170;48;5;235m▒\033[38;5;95;48;5;235m▓\033[38;5;208;48;5;94m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;222m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;94m▒\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;172m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;137m▒\033[38;5;209;48;5;234m▓\033[38;5;204;48;5;235m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;220;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;221m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;208;48;5;94m▒\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m░\033[38;5;173;48;5;235m▓\033[38;5;61;48;5;235m▒\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;161;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m \033[38;5;137;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;137;48;5;237m▒\033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;166;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;61;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;180;48;5;58m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;94;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m░\033[38;5;204;48;5;234m▓\033[38;5;95;48;5;235m▓\033[38;5;172;48;5;137m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;208;48;5;94m░\033[38;5;209;48;5;235m▓\033[38;5;48;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;168;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;236m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;136;48;5;229m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;94m▒\033[38;5;204;48;5;234m▓\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;130m░\033[38;5;209;48;5;235m▓\033[38;5;133;48;5;235m▓\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;78;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;208;48;5;94m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;221m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;229m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;137m▒\033[38;5;209;48;5;234m▓\033[38;5;166;48;5;236m▒\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m▒\033[38;5;204;48;5;234m▓\033[38;5;104;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;161;48;5;235m▒\033[38;5;173;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;130;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;173m▒\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;173m▒\033[38;5;95;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;204;48;5;235m░\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;234m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;208;48;5;130m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;209;48;5;234m▒\033[38;5;133;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;166;48;5;237m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;214;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;208;48;5;130m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;202;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;94m▒\033[38;5;202;48;5;236m▓\033[38;5;95;48;5;234m▓\033[38;5;95;48;5;234m▓\033[38;5;166;48;5;236m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;180;48;5;58m▒\033[38;5;209;48;5;235m▓\033[38;5;126;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;133;48;5;235m▓\033[38;5;95;48;5;234m▓\033[38;5;130;48;5;95m▒\033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;173m░\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;94m▒\033[38;5;166;48;5;237m▒\033[38;5;166;48;5;237m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;136;48;5;229m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;223m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;179m░\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;101;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;179m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;136;48;5;229m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;58m▒\033[38;5;209;48;5;235m▓\033[38;5;98;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;168;48;5;235m▒\033[38;5;95;48;5;235m▓\033[38;5;130;48;5;58m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;137m▒\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;234m▒\033[38;5;69;48;5;235m▒\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;172m░\033[38;5;130;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;173;48;5;235m▓\033[38;5;172;48;5;179m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;173;48;5;235m▓\033[38;5;104;48;5;235m▒\033[38;5;167;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;234m▒\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;236m▓\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;237m▒\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;220;48;5;230m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;130m▒\033[38;5;209;48;5;235m▓\033[38;5;47;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;98;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m░\033[38;5;130;48;5;214m░\033[38;5;137;48;5;237m▒\033[38;5;204;48;5;234m▓\033[38;5;130;48;5;173m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;94;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m░\033[38;5;209;48;5;235m▓\033[38;5;129;48;5;235m▓\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;202;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;208;48;5;94m▒\033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;208;48;5;94m░\033[38;5;204;48;5;234m▓\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;229m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;166;48;5;236m▒\033[38;5;209;48;5;235m▓\033[38;5;167;48;5;233m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;84;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;130;48;5;130m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;166m░\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;236m▓\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;208;48;5;94m░\033[38;5;95;48;5;235m▓\033[38;5;42;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;214;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;208;48;5;58m▒\033[38;5;95;48;5;235m▓\033[38;5;208;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;173;48;5;235m▓\033[38;5;61;48;5;235m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;69;48;5;235m▒\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;214m░\033[38;5;172;48;5;214m \033[38;5;172;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;172m░\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;236m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;223m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;166;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;190;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;234m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;208;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;208;48;5;94m░\033[38;5;204;48;5;234m▓\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;208;48;5;94m░\033[38;5;209;48;5;235m▓\033[38;5;197;48;5;235m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;98;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;180;48;5;58m▒\033[38;5;95;48;5;234m▓\033[38;5;208;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;94;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;173m▒\033[38;5;173;48;5;235m▓\033[38;5;104;48;5;235m▒\033[38;5;167;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;175;48;5;235m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;58m▒\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;137;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;222m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;137;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;129;48;5;235m░\033[38;5;173;48;5;238m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;252m▓\033[38;5;209;48;5;233m▒\033[38;5;209;48;5;234m▒\033[38;5;166;48;5;188m▓\033[38;5;209;48;5;237m▓\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;173m░\033[38;5;130;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;214m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;214m░\033[38;5;130;48;5;214m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;230m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;94m▒\033[38;5;95;48;5;235m▓\033[38;5;78;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;41;48;5;237m▒\033[38;5;173;48;5;234m▓\033[38;5;202;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;223;48;5;224m░\033[38;5;173;48;5;237m▓\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;173m░\033[38;5;130;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;94;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;130m░\033[38;5;209;48;5;235m▓\033[38;5;175;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;234m▒\033[38;5;55;48;5;235m░\033[38;5;173;48;5;237m▓\033[38;5;166;48;5;253m▒\033[38;5;223;48;5;230m \033[38;5;180;48;5;224m▒\033[38;5;180;48;5;224m▒\033[38;5;166;48;5;224m░\033[38;5;173;48;5;238m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;180;48;5;237m▒\033[38;5;46;48;5;235m░\033[38;5;209;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;72;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;234m▓\033[38;5;173;48;5;234m▓\033[38;5;173;48;5;234m▓\033[38;5;173;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;172;48;5;172m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;62;48;5;208m░\033[38;5;204;48;5;208m░\033[38;5;48;48;5;209m░\033[38;5;121;48;5;209m░\033[38;5;42;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;1;48;5;232m░\033[0m░\033[0m░\033[38;5;209;48;5;236m▓\033[0m \033[0m \033[0m \033[38;5;131;48;5;236m▒\033[38;5;180;48;5;236m▒\033[38;5;179;48;5;52m▒\033[38;5;29;48;5;222m░\033[38;5;41;48;5;209m░\033[38;5;35;48;5;209m░\033[38;5;163;48;5;208m \033[38;5;169;48;5;208m▒\033[38;5;62;48;5;208m▒\033[38;5;81;48;5;208m▒\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;51;48;5;231m░\033[38;5;51;48;5;231m░\033[38;5;51;48;5;231m░\033[38;5;51;48;5;231m░\033[38;5;82;48;5;215m░\033[38;5;80;48;5;215m▒\033[38;5;220;48;5;221m░\033[38;5;122;48;5;215m░\033[38;5;48;48;5;208m░\033[38;5;41;48;5;209m░\033[38;5;43;48;5;223m░\033[38;5;179;48;5;236m▒\033[38;5;130;48;5;52m▒\033[38;5;173;48;5;237m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;173;48;5;240m▓\033[38;5;73;48;5;249m▓\033[38;5;73;48;5;249m▓\033[38;5;73;48;5;249m▓\033[38;5;73;48;5;249m▓\033[38;5;73;48;5;249m▓\033[38;5;73;48;5;249m▓\033[38;5;73;48;5;249m▓\033[38;5;73;48;5;249m▓\033[38;5;73;48;5;249m▓\033[38;5;73;48;5;249m▓\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m");
end
endtask

task FAIL;
begin
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;167;48;5;234m▒\033[38;5;202;48;5;234m▓\033[38;5;48;48;5;236m▓\033[38;5;161;48;5;235m▒\033[38;5;98;48;5;235m▓\033[38;5;69;48;5;235m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;69;48;5;235m▒\033[38;5;98;48;5;235m▓\033[38;5;169;48;5;235m▒\033[38;5;35;48;5;236m▓\033[38;5;202;48;5;234m▓\033[38;5;209;48;5;234m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;209;48;5;235m▒\033[38;5;208;48;5;236m▓\033[38;5;202;48;5;236m▓\033[38;5;209;48;5;235m▒\033[38;5;52;48;5;232m░\033[38;5;52;48;5;232m░\033[38;5;1;48;5;232m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;52;48;5;232m░\033[38;5;190;48;5;236m▓\033[38;5;168;48;5;235m▒\033[38;5;69;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;236m▒\033[38;5;208;48;5;238m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;173m▒\033[38;5;208;48;5;130m░\033[38;5;208;48;5;94m░\033[38;5;180;48;5;237m▒\033[38;5;166;48;5;236m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;69;48;5;235m▒\033[38;5;161;48;5;235m▒\033[38;5;112;48;5;236m▓\033[38;5;52;48;5;232m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;1;48;5;232m░\033[38;5;52;48;5;232m░\033[38;5;52;48;5;232m░\033[38;5;209;48;5;234m▒\033[38;5;202;48;5;236m▓\033[38;5;137;48;5;236m▓\033[38;5;209;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;206;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;137;48;5;237m▒\033[38;5;166;48;5;237m▒\033[38;5;202;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;129;48;5;235m▓\033[38;5;35;48;5;236m▓\033[38;5;166;48;5;236m▓\033[38;5;167;48;5;233m░\033[38;5;1;48;5;232m░\033[38;5;179;48;5;236m▓\033[38;5;133;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;208;48;5;238m▒\033[38;5;130;48;5;136m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;137m▒\033[38;5;130;48;5;58m▒\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;99;48;5;235m▒\033[38;5;221;48;5;236m▓\033[38;5;1;48;5;232m░\033[0m \033[38;5;173;48;5;236m▓\033[38;5;35;48;5;236m▓\033[38;5;133;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;236m▓\033[38;5;166;48;5;237m▒\033[38;5;137;48;5;237m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;104;48;5;235m▒\033[0m░\033[0m \033[0m \033[38;5;243;48;5;242m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;236m▒\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;240m▓\033[38;5;204;48;5;175m▒\033[38;5;204;48;5;95m▓\033[38;5;202;48;5;236m▓\033[38;5;172;48;5;173m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;179m░\033[38;5;172;48;5;137m▒\033[38;5;180;48;5;238m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;173m░\033[38;5;130;48;5;58m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;166;48;5;237m▒\033[38;5;172;48;5;137m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;173m░\033[38;5;166;48;5;236m▒\033[38;5;204;48;5;240m▓\033[38;5;204;48;5;174m▒\033[38;5;204;48;5;95m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;130;48;5;236m▓\033[38;5;173;48;5;234m▓\033[38;5;204;48;5;95m▓\033[38;5;168;48;5;211m░\033[38;5;204;48;5;175m░\033[38;5;204;48;5;211m░\033[38;5;204;48;5;132m▓\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;137m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;173m░\033[38;5;180;48;5;238m▒\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;137;48;5;237m▒\033[38;5;172;48;5;137m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;214m \033[38;5;172;48;5;214m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;173m▒\033[38;5;180;48;5;238m▒\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;137;48;5;237m▒\033[38;5;172;48;5;173m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;137m▒\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;131m▓\033[38;5;204;48;5;175m░\033[38;5;204;48;5;175m░\033[38;5;204;48;5;211m░\033[38;5;168;48;5;132m▓\033[38;5;173;48;5;234m▓\033[38;5;190;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;76;48;5;236m▓\033[38;5;173;48;5;234m▓\033[38;5;197;48;5;132m▓\033[38;5;218;48;5;218m \033[38;5;161;48;5;218m \033[38;5;168;48;5;211m░\033[38;5;204;48;5;211m░\033[38;5;204;48;5;211m░\033[38;5;204;48;5;132m▓\033[38;5;202;48;5;236m▓\033[38;5;130;48;5;94m▒\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;236m▒\033[38;5;172;48;5;179m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;180;48;5;238m▒\033[38;5;95;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;180;48;5;238m▒\033[38;5;166;48;5;237m▓\033[38;5;204;48;5;131m▓\033[38;5;204;48;5;211m░\033[38;5;204;48;5;175m░\033[38;5;204;48;5;175m░\033[38;5;197;48;5;211m░\033[38;5;218;48;5;218m \033[38;5;168;48;5;174m▒\033[38;5;173;48;5;234m▓\033[38;5;48;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;78;48;5;236m▓\033[38;5;173;48;5;234m▓\033[38;5;197;48;5;132m▓\033[38;5;218;48;5;218m \033[38;5;218;48;5;218m \033[38;5;218;48;5;218m \033[38;5;161;48;5;218m \033[38;5;204;48;5;174m▒\033[38;5;138;48;5;238m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;137m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;137m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;131m▒\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;173m▒\033[38;5;166;48;5;236m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;236m▓\033[38;5;204;48;5;132m▓\033[38;5;197;48;5;211m \033[38;5;161;48;5;218m \033[38;5;218;48;5;218m \033[38;5;218;48;5;218m \033[38;5;168;48;5;174m▒\033[38;5;173;48;5;234m▓\033[38;5;35;48;5;235m▒\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;78;48;5;236m▓\033[38;5;173;48;5;234m▓\033[38;5;197;48;5;132m▓\033[38;5;218;48;5;218m \033[38;5;218;48;5;218m \033[38;5;197;48;5;211m░\033[38;5;204;48;5;239m▓\033[38;5;173;48;5;235m▓\033[38;5;166;48;5;236m▓\033[38;5;172;48;5;173m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;94m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;131m▒\033[38;5;130;48;5;58m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;208;48;5;238m▒\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;236m▓\033[38;5;197;48;5;175m▒\033[38;5;218;48;5;218m \033[38;5;218;48;5;218m \033[38;5;168;48;5;174m▒\033[38;5;173;48;5;234m▓\033[38;5;35;48;5;235m▒\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;78;48;5;236m▓\033[38;5;173;48;5;234m▓\033[38;5;197;48;5;132m▓\033[38;5;198;48;5;218m \033[38;5;168;48;5;96m▓\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;173m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;166;48;5;236m▓\033[38;5;130;48;5;131m▒\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;137m▒\033[38;5;173;48;5;235m▓\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;166;48;5;236m▒\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;239m▓\033[38;5;161;48;5;218m \033[38;5;168;48;5;174m▒\033[38;5;173;48;5;234m▓\033[38;5;35;48;5;235m▒\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;78;48;5;236m▓\033[38;5;173;48;5;234m▓\033[38;5;204;48;5;132m▓\033[38;5;204;48;5;237m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;58m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;172;48;5;137m▒\033[38;5;166;48;5;237m▒\033[38;5;208;48;5;238m▒\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;94;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m▒\033[38;5;208;48;5;58m▒\033[38;5;166;48;5;237m▒\033[38;5;130;48;5;95m▒\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;137m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;236m▓\033[38;5;204;48;5;95m▓\033[38;5;173;48;5;235m▓\033[38;5;42;48;5;235m▒\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;191;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;137m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;94m▒\033[38;5;166;48;5;236m▒\033[38;5;180;48;5;238m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;94m▒\033[38;5;180;48;5;238m▒\033[38;5;166;48;5;236m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;173m░\033[38;5;202;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;84;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;130;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;173m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;230;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;202;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;35;48;5;235m▓\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;234m▒\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;172;48;5;173m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;137m▒\033[38;5;208;48;5;238m▒\033[38;5;202;48;5;59m▓\033[38;5;173;48;5;240m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;242m▓\033[38;5;166;48;5;224m▒\033[38;5;166;48;5;187m▓\033[38;5;202;48;5;243m▓\033[38;5;180;48;5;238m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;58m▒\033[38;5;202;48;5;242m▓\033[38;5;166;48;5;187m▓\033[38;5;166;48;5;224m▒\033[38;5;202;48;5;244m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;239m▓\033[38;5;166;48;5;59m▓\033[38;5;166;48;5;238m▓\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;82;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;99;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;208;48;5;130m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;166;48;5;238m▒\033[38;5;202;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;245m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;255;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;249m▓\033[38;5;166;48;5;238m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;223m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;180;48;5;238m▒\033[38;5;209;48;5;247m▓\033[38;5;231;48;5;231m▓\033[38;5;137;48;5;255m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;243m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;180;48;5;254m▒\033[38;5;166;48;5;238m▓\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;208;48;5;130m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;65;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;236m▒\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;208;48;5;239m▒\033[38;5;173;48;5;242m▓\033[38;5;209;48;5;249m▓\033[38;5;209;48;5;247m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;202;48;5;236m▓\033[38;5;208;48;5;238m▒\033[38;5;130;48;5;94m▒\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;131m▒\033[38;5;208;48;5;238m▒\033[38;5;166;48;5;236m▓\033[38;5;166;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;173;48;5;246m▓\033[38;5;166;48;5;7m▓\033[38;5;202;48;5;242m▓\033[38;5;137;48;5;238m▒\033[38;5;172;48;5;179m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;180;48;5;58m▒\033[38;5;209;48;5;235m▓\033[38;5;197;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;99;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;208;48;5;130m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;94;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;255m▓\033[38;5;173;48;5;251m▓\033[38;5;173;48;5;248m▓\033[38;5;166;48;5;247m▓\033[38;5;173;48;5;250m▓\033[38;5;95;48;5;255m▓\033[38;5;209;48;5;253m▓\033[38;5;209;48;5;145m▓\033[38;5;173;48;5;248m▓\033[38;5;202;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;224;48;5;231m \033[38;5;209;48;5;188m▓\033[38;5;209;48;5;249m▓\033[38;5;209;48;5;249m▓\033[38;5;209;48;5;251m▓\033[38;5;173;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;223m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;232m░\033[38;5;173;48;5;235m▓\033[38;5;202;48;5;236m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;136;48;5;229m \033[38;5;231;48;5;231m▓\033[38;5;173;48;5;254m▓\033[38;5;173;48;5;240m▓\033[38;5;173;48;5;242m▓\033[38;5;209;48;5;251m▓\033[38;5;216;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;255;48;5;255m▓\033[38;5;209;48;5;237m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;173;48;5;242m▓\033[38;5;179;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;137;48;5;231m▓\033[38;5;209;48;5;251m▓\033[38;5;209;48;5;240m▓\033[38;5;209;48;5;59m▓\033[38;5;138;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;94;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;166;48;5;58m▒\033[38;5;209;48;5;235m▓\033[38;5;35;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;113;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;180;48;5;237m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;246m▓\033[38;5;209;48;5;241m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;240m▓\033[38;5;253;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;137;48;5;231m▓\033[38;5;173;48;5;237m▓\033[38;5;173;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;130m▒\033[38;5;209;48;5;235m▓\033[38;5;133;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;84;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;222m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;239m▓\033[38;5;209;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;241m▓\033[38;5;209;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;166;48;5;7m▓\033[38;5;173;48;5;241m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;249m▓\033[38;5;166;48;5;254m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;230m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;214m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m▒\033[38;5;173;48;5;235m▓\033[38;5;104;48;5;235m▒\033[38;5;167;48;5;233m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;113;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;180;48;5;238m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;178;48;5;229m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;59m▓\033[38;5;209;48;5;247m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;130;48;5;255m \033[38;5;173;48;5;246m▓\033[38;5;173;48;5;235m▓\033[38;5;202;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;247m▓\033[38;5;209;48;5;243m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;255m▓\033[38;5;173;48;5;235m▓\033[38;5;166;48;5;188m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;137m▒\033[38;5;209;48;5;235m▓\033[38;5;69;48;5;235m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;173;48;5;235m▓\033[38;5;166;48;5;236m▓\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;239m▓\033[38;5;173;48;5;241m▓\033[38;5;180;48;5;224m▒\033[38;5;166;48;5;224m░\033[38;5;166;48;5;255m \033[38;5;166;48;5;230m \033[38;5;166;48;5;224m░\033[38;5;166;48;5;224m░\033[38;5;166;48;5;224m░\033[38;5;166;48;5;253m▒\033[38;5;173;48;5;239m▓\033[38;5;204;48;5;95m▓\033[38;5;204;48;5;211m░\033[38;5;204;48;5;95m▓\033[38;5;173;48;5;236m▓\033[38;5;166;48;5;187m▓\033[38;5;166;48;5;224m░\033[38;5;166;48;5;224m░\033[38;5;166;48;5;224m░\033[38;5;166;48;5;230m \033[38;5;166;48;5;255m \033[38;5;166;48;5;224m░\033[38;5;166;48;5;224m░\033[38;5;166;48;5;144m▓\033[38;5;209;48;5;237m▓\033[38;5;95;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;238m▓\033[38;5;166;48;5;248m▓\033[38;5;222;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;178;48;5;230m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;130m▒\033[38;5;209;48;5;235m▓\033[38;5;98;48;5;235m▓\033[38;5;209;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;99;48;5;235m░\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;136;48;5;229m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;202;48;5;138m▓\033[38;5;173;48;5;239m▓\033[38;5;209;48;5;237m▓\033[38;5;209;48;5;237m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;237m▓\033[38;5;209;48;5;237m▓\033[38;5;204;48;5;95m▓\033[38;5;168;48;5;211m░\033[38;5;161;48;5;218m \033[38;5;161;48;5;218m \033[38;5;197;48;5;211m░\033[38;5;168;48;5;175m▒\033[38;5;209;48;5;236m▓\033[38;5;173;48;5;239m▓\033[38;5;209;48;5;237m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;236m▓\033[38;5;173;48;5;236m▓\033[38;5;173;48;5;238m▓\033[38;5;202;48;5;243m▓\033[38;5;166;48;5;252m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;255m▓\033[38;5;173;48;5;236m▓\033[38;5;166;48;5;252m▒\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;58m▒\033[38;5;209;48;5;235m▓\033[38;5;49;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m░\033[0m \033[38;5;42;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;208;48;5;58m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;221;48;5;223m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;216;48;5;231m \033[38;5;181;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;237m▓\033[38;5;197;48;5;211m░\033[38;5;218;48;5;218m \033[38;5;218;48;5;218m \033[38;5;218;48;5;218m \033[38;5;168;48;5;132m▓\033[38;5;209;48;5;242m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;202;48;5;254m▓\033[38;5;221;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;172m░\033[38;5;202;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;172m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;246m▓\033[38;5;173;48;5;241m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;236m▓\033[38;5;173;48;5;238m▓\033[38;5;173;48;5;237m▓\033[38;5;209;48;5;234m▓\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;188m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;137;48;5;231m▓\033[38;5;173;48;5;237m▓\033[38;5;168;48;5;132m▓\033[38;5;197;48;5;175m▒\033[38;5;204;48;5;95m▓\033[38;5;209;48;5;240m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;221;48;5;223m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;180;48;5;94m░\033[38;5;209;48;5;235m▓\033[38;5;91;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;29;48;5;235m▒\033[38;5;173;48;5;235m▓\033[38;5;180;48;5;58m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;94;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;242m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;102m▓\033[38;5;173;48;5;243m▓\033[38;5;209;48;5;239m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;243m▓\033[38;5;209;48;5;234m▓\033[38;5;166;48;5;245m▓\033[38;5;166;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;229m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;214m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;222m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;137;48;5;254m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;239m▓\033[38;5;209;48;5;188m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;249m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;246m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;238m▓\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;145m▓\033[38;5;172;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;222m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;208;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;202;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;65;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;202;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;230;48;5;230m \033[38;5;173;48;5;249m▓\033[38;5;209;48;5;253m▓\033[38;5;209;48;5;243m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;236m▓\033[38;5;166;48;5;242m▓\033[38;5;208;48;5;255m \033[38;5;231;48;5;231m▓\033[38;5;209;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;166;48;5;224m░\033[38;5;202;48;5;236m▓\033[38;5;173;48;5;237m▓\033[38;5;166;48;5;188m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;229m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;202;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;72;48;5;235m▓\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;137;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;208;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;95;48;5;255m▓\033[38;5;137;48;5;254m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;244m▓\033[38;5;172;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;243m▓\033[38;5;209;48;5;234m▓\033[38;5;202;48;5;246m▓\033[38;5;223;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;136;48;5;229m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;137m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;84;48;5;236m▓\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;136;48;5;229m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;238m▓\033[38;5;209;48;5;242m▓\033[38;5;209;48;5;253m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;202;48;5;247m▓\033[38;5;209;48;5;234m▓\033[38;5;173;48;5;243m▓\033[38;5;166;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;94m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;133;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;236m▓\033[38;5;130;48;5;173m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;94;48;5;223m \033[38;5;209;48;5;239m▓\033[38;5;209;48;5;239m▓\033[38;5;178;48;5;230m \033[38;5;136;48;5;229m \033[38;5;94;48;5;222m \033[38;5;94;48;5;222m \033[38;5;222;48;5;222m \033[38;5;222;48;5;222m \033[38;5;94;48;5;222m \033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;173;48;5;245m▓\033[38;5;209;48;5;234m▓\033[38;5;202;48;5;245m▓\033[38;5;166;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;137m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;35;48;5;235m▒\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;173;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;202;48;5;236m▓\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;180;48;5;238m▒\033[38;5;166;48;5;236m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;222m \033[38;5;209;48;5;241m▓\033[38;5;209;48;5;234m▓\033[38;5;166;48;5;145m▓\033[38;5;223;48;5;230m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;214;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;94m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;168;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;232m░\033[38;5;133;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;173m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;94m▒\033[38;5;95;48;5;234m▓\033[38;5;172;48;5;179m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;137;48;5;237m▒\033[38;5;209;48;5;236m▓\033[38;5;166;48;5;187m▓\033[38;5;208;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;230m \033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;179m░\033[38;5;130;48;5;94m▒\033[38;5;202;48;5;236m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;65;48;5;235m▓\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;119;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;173m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m▒\033[38;5;209;48;5;235m▓\033[38;5;180;48;5;94m▒\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;239m▓\033[38;5;166;48;5;224m▒\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m▒\033[38;5;208;48;5;58m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;191;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;48;48;5;235m▓\033[38;5;104;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;69;48;5;235m▒\033[38;5;98;48;5;235m▓\033[38;5;79;48;5;235m▒\033[38;5;209;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;168;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;131m▒\033[38;5;130;48;5;173m░\033[38;5;130;48;5;94m▒\033[38;5;166;48;5;236m▒\033[38;5;95;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;208;48;5;238m▒\033[38;5;202;48;5;236m▒\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;94m░\033[38;5;209;48;5;234m▓\033[38;5;202;48;5;245m▓\033[38;5;166;48;5;224m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m░\033[38;5;130;48;5;94m▒\033[38;5;209;48;5;235m▓\033[38;5;204;48;5;234m▓\033[38;5;95;48;5;235m▓\033[38;5;166;48;5;237m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;166;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;221;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;72;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;236m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;137m▒\033[38;5;172;48;5;173m▒\033[38;5;172;48;5;179m░\033[38;5;172;48;5;179m░\033[38;5;172;48;5;179m░\033[38;5;172;48;5;173m▒\033[38;5;130;48;5;136m▒\033[38;5;208;48;5;94m░\033[38;5;166;48;5;237m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;168;48;5;235m▒\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;101;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;208;48;5;58m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;94m▒\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;173m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;166;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;246m▓\033[38;5;166;48;5;251m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;230;48;5;231m \033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m▒\033[38;5;173;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;35;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;137;48;5;237m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;130m░\033[38;5;166;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;235m▒\033[38;5;69;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;173m░\033[38;5;166;48;5;236m▒\033[38;5;180;48;5;238m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;172m░\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;238m▓\033[38;5;173;48;5;244m▓\033[38;5;173;48;5;239m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;239m▓\033[38;5;137;48;5;255m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;188m▓\033[38;5;202;48;5;245m▓\033[38;5;209;48;5;240m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;234m▓\033[38;5;204;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;166;48;5;237m▒\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;136m▒\033[38;5;209;48;5;235m▓\033[38;5;61;48;5;235m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;1;48;5;232m░\033[38;5;169;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;137;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;99;48;5;235m▒\033[38;5;52;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[38;5;119;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;208;48;5;58m▒\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;130m▒\033[38;5;95;48;5;235m▓\033[38;5;172;48;5;137m▒\033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;208;48;5;58m▒\033[38;5;209;48;5;234m▓\033[38;5;166;48;5;249m▓\033[38;5;166;48;5;224m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;173;48;5;242m▓\033[38;5;209;48;5;234m▓\033[38;5;173;48;5;236m▓\033[38;5;173;48;5;239m▓\033[38;5;209;48;5;240m▓\033[38;5;209;48;5;238m▓\033[38;5;173;48;5;237m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;234m▓\033[38;5;209;48;5;234m▓\033[38;5;202;48;5;236m▓\033[38;5;208;48;5;58m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;179m░\033[38;5;137;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;172;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;236m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;173m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;172m░\033[38;5;208;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;166;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;79;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[38;5;98;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;208;48;5;238m▒\033[38;5;202;48;5;235m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;136m░\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;239m▓\033[38;5;166;48;5;224m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;209;48;5;244m▓\033[38;5;202;48;5;247m▓\033[38;5;172;48;5;179m░\033[38;5;172;48;5;179m░\033[38;5;172;48;5;179m░\033[38;5;130;48;5;173m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;130;48;5;137m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;167;48;5;233m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;41;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;166;48;5;237m▒\033[38;5;208;48;5;94m░\033[38;5;208;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;94m▒\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;119;48;5;235m▓\033[38;5;209;48;5;236m▒\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;236m▒\033[38;5;130;48;5;172m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;179m░\033[38;5;202;48;5;236m▓\033[38;5;180;48;5;237m▒\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;208;48;5;94m░\033[38;5;95;48;5;235m▓\033[38;5;166;48;5;138m▓\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;222;48;5;221m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;180;48;5;58m▒\033[38;5;209;48;5;235m▓\033[38;5;65;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[0m░\033[38;5;209;48;5;236m▒\033[38;5;209;48;5;236m▒\033[38;5;208;48;5;236m▓\033[38;5;42;48;5;235m▒\033[38;5;104;48;5;235m▒\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;166;48;5;236m▒\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;208;48;5;94m░\033[38;5;130;48;5;172m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;173m▒\033[38;5;138;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;172m░\033[38;5;180;48;5;58m▒\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;145m▓\033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;94;48;5;223m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;172m░\033[38;5;130;48;5;130m░\033[38;5;95;48;5;235m▓\033[38;5;69;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;233m░\033[38;5;129;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;236m▓\033[38;5;130;48;5;173m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;173m▒\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;94m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;215m░\033[38;5;130;48;5;94m▒\033[38;5;95;48;5;235m▓\033[38;5;202;48;5;243m▓\033[38;5;166;48;5;188m▒\033[38;5;166;48;5;224m░\033[38;5;166;48;5;255m \033[38;5;223;48;5;255m \033[38;5;178;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;214;48;5;222m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;166;48;5;236m▒\033[38;5;173;48;5;235m▓\033[38;5;101;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;78;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;208;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;173m░\033[38;5;95;48;5;235m▓\033[38;5;180;48;5;237m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;222;48;5;215m \033[38;5;172;48;5;215m░\033[38;5;202;48;5;235m▓\033[38;5;208;48;5;238m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;179m░\033[38;5;130;48;5;180m▒\033[38;5;202;48;5;245m▓\033[38;5;209;48;5;236m▓\033[38;5;209;48;5;234m▓\033[38;5;173;48;5;239m▓\033[38;5;202;48;5;247m▓\033[38;5;130;48;5;180m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;173m░\033[38;5;130;48;5;173m▒\033[38;5;130;48;5;137m▒\033[38;5;208;48;5;58m▒\033[38;5;173;48;5;236m▓\033[38;5;95;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;208;48;5;58m▒\033[38;5;172;48;5;173m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;208;48;5;94m░\033[38;5;209;48;5;235m▓\033[38;5;197;48;5;235m▒\033[38;5;88;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;84;48;5;236m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;130m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;130m▒\033[38;5;204;48;5;234m▓\033[38;5;208;48;5;94m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;214m \033[38;5;130;48;5;94m▒\033[38;5;130;48;5;58m▒\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;214;48;5;221m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;223;48;5;255m \033[38;5;166;48;5;224m░\033[38;5;166;48;5;248m▓\033[38;5;209;48;5;239m▓\033[38;5;209;48;5;235m▓\033[38;5;209;48;5;234m▓\033[38;5;204;48;5;234m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;236m▓\033[38;5;166;48;5;236m▒\033[38;5;166;48;5;237m▒\033[38;5;166;48;5;237m▒\033[38;5;180;48;5;58m▒\033[38;5;180;48;5;58m▒\033[38;5;180;48;5;58m▒\033[38;5;137;48;5;237m▒\033[38;5;166;48;5;236m▒\033[38;5;166;48;5;236m▓\033[38;5;173;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;95;48;5;235m▓\033[38;5;204;48;5;234m▓\033[38;5;204;48;5;234m▓\033[38;5;95;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;166;48;5;236m▒\033[38;5;130;48;5;94m▒\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;179m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;130;48;5;130m░\033[38;5;209;48;5;235m▓\033[38;5;69;48;5;235m▒\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;130;48;5;234m▓\033[38;5;209;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;130;48;5;130m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;137;48;5;237m▒\033[38;5;95;48;5;235m▓\033[38;5;130;48;5;130m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m \033[38;5;222;48;5;215m \033[38;5;130;48;5;215m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;216;48;5;203m \033[38;5;220;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;209;48;5;217m▒\033[38;5;166;48;5;252m▒\033[38;5;166;48;5;187m▓\033[38;5;166;48;5;181m▓\033[38;5;166;48;5;181m▓\033[38;5;166;48;5;249m▓\033[38;5;166;48;5;145m▓\033[38;5;202;48;5;145m▓\033[38;5;204;48;5;203m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;203;48;5;209m░\033[38;5;166;48;5;224m▒\033[38;5;166;48;5;224m▒\033[38;5;166;48;5;224m░\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;209;48;5;202m░\033[38;5;172;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;202;48;5;236m▓\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;234m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;202;48;5;235m▓\033[38;5;173;48;5;235m▓\033[38;5;209;48;5;235m▓\033[38;5;130;48;5;137m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;179m░\033[38;5;209;48;5;235m▓\033[38;5;202;48;5;236m▒\033[38;5;130;48;5;172m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;215;48;5;208m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;196;48;5;196m \033[38;5;196;48;5;196m \033[38;5;196;48;5;196m \033[38;5;196;48;5;196m \033[38;5;196;48;5;196m \033[38;5;196;48;5;196m \033[38;5;216;48;5;209m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;217m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;203m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;210m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;209;48;5;202m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;130;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;172m░\033[38;5;180;48;5;237m▒\033[38;5;209;48;5;235m▓\033[38;5;84;48;5;236m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;52;48;5;232m░\033[38;5;61;48;5;235m▒\033[38;5;209;48;5;235m▓\033[38;5;208;48;5;238m▒\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;215m░\033[38;5;130;48;5;137m▒\033[38;5;204;48;5;235m▓\033[38;5;208;48;5;238m▒\033[38;5;172;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;166;48;5;208m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;178;48;5;230m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;203m \033[38;5;204;48;5;210m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;217m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;210m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;209;48;5;202m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;214m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;94m▒\033[38;5;209;48;5;235m▓\033[38;5;35;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;113;48;5;236m▓\033[38;5;104;48;5;235m▒\033[38;5;209;48;5;237m░\033[38;5;79;48;5;137m▓\033[38;5;202;48;5;239m▓\033[0m░\033[38;5;52;48;5;232m░\033[38;5;1;48;5;232m░\033[38;5;43;48;5;186m░\033[38;5;64;48;5;215m░\033[38;5;222;48;5;215m░\033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;166;48;5;208m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;221m \033[38;5;230;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;231m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;210m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;209;48;5;202m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;172;48;5;215m \033[38;5;130;48;5;131m▒\033[38;5;209;48;5;235m▓\033[38;5;42;48;5;235m▒\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;131;48;5;237m▒\033[38;5;42;48;5;137m▒\033[38;5;35;48;5;137m▒\033[38;5;42;48;5;137m▒\033[38;5;36;48;5;221m░\033[38;5;45;48;5;215m░\033[38;5;172;48;5;215m░\033[38;5;130;48;5;214m \033[38;5;215;48;5;208m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;204m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;217m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;224m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;203m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;210m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;209;48;5;202m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;208m░\033[38;5;130;48;5;214m░\033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m░\033[38;5;43;48;5;222m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m░\033[38;5;216;48;5;233m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;255m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;203m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;210m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;210m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;209;48;5;202m \033[38;5;130;48;5;214m░\033[38;5;130;48;5;214m \033[38;5;172;48;5;215m \033[38;5;172;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m \033[38;5;222;48;5;215m░\033[38;5;45;48;5;215m░\033[38;5;86;48;5;215m░\033[38;5;29;48;5;221m░\033[38;5;29;48;5;215m░\033[38;5;86;48;5;102m▓\033[0m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;232m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;167;48;5;234m▒\033[38;5;108;48;5;95m▓\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;231m░\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;210m \033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;231;48;5;231m▓\033[38;5;204;48;5;203m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;84;48;5;202m░\033[38;5;86;48;5;215m░\033[38;5;36;48;5;222m░\033[38;5;50;48;5;223m░\033[38;5;178;48;5;237m▓\033[38;5;209;48;5;239m▓\033[38;5;95;48;5;240m▓\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;232m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;137;48;5;196m▓\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;119;48;5;88m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m░\033[38;5;1;48;5;232m░\033[0m \033[0m \033[38;5;35;48;5;196m▓\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;46;48;5;196m░\033[0m \033[0m \033[0m \033[38;5;204;48;5;196m▒\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;50;48;5;196m▒\033[38;5;46;48;5;196m░\033[38;5;46;48;5;196m░\033[38;5;46;48;5;196m░\033[38;5;46;48;5;196m░\033[38;5;46;48;5;196m░\033[38;5;46;48;5;196m░\033[38;5;64;48;5;52m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;209;48;5;232m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;82;48;5;52m░\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;130;48;5;52m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[38;5;47;48;5;196m▒\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m░\033[0m \033[0m \033[38;5;35;48;5;196m▓\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;46;48;5;196m░\033[0m \033[0m \033[0m \033[38;5;204;48;5;196m▒\033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;204;48;5;196m \033[38;5;76;48;5;52m░\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m \033[0m");
$display("\033[0m");
end
endtask

endmodule
